magic
tech sky130A
magscale 1 2
timestamp 1647671105
<< obsli1 >>
rect 1104 2159 65412 66385
<< obsm1 >>
rect 658 2128 65766 66416
<< metal2 >>
rect 634 67943 746 68743
rect 1922 67943 2034 68743
rect 3210 67943 3322 68743
rect 4498 67943 4610 68743
rect 5786 67943 5898 68743
rect 7074 67943 7186 68743
rect 8362 67943 8474 68743
rect 9650 67943 9762 68743
rect 10294 67943 10406 68743
rect 11582 67943 11694 68743
rect 12870 67943 12982 68743
rect 14158 67943 14270 68743
rect 15446 67943 15558 68743
rect 16734 67943 16846 68743
rect 18022 67943 18134 68743
rect 19310 67943 19422 68743
rect 20598 67943 20710 68743
rect 21886 67943 21998 68743
rect 23174 67943 23286 68743
rect 24462 67943 24574 68743
rect 25750 67943 25862 68743
rect 27038 67943 27150 68743
rect 28326 67943 28438 68743
rect 28970 67943 29082 68743
rect 30258 67943 30370 68743
rect 31546 67943 31658 68743
rect 32834 67943 32946 68743
rect 34122 67943 34234 68743
rect 35410 67943 35522 68743
rect 36698 67943 36810 68743
rect 37986 67943 38098 68743
rect 39274 67943 39386 68743
rect 40562 67943 40674 68743
rect 41850 67943 41962 68743
rect 43138 67943 43250 68743
rect 44426 67943 44538 68743
rect 45714 67943 45826 68743
rect 47002 67943 47114 68743
rect 47646 67943 47758 68743
rect 48934 67943 49046 68743
rect 50222 67943 50334 68743
rect 51510 67943 51622 68743
rect 52798 67943 52910 68743
rect 54086 67943 54198 68743
rect 55374 67943 55486 68743
rect 56662 67943 56774 68743
rect 57950 67943 58062 68743
rect 59238 67943 59350 68743
rect 60526 67943 60638 68743
rect 61814 67943 61926 68743
rect 63102 67943 63214 68743
rect 64390 67943 64502 68743
rect 65678 67943 65790 68743
rect 66322 67943 66434 68743
rect -10 0 102 800
rect 634 0 746 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 4498 0 4610 800
rect 5786 0 5898 800
rect 7074 0 7186 800
rect 8362 0 8474 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 12226 0 12338 800
rect 13514 0 13626 800
rect 14802 0 14914 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 21886 0 21998 800
rect 23174 0 23286 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 34766 0 34878 800
rect 36054 0 36166 800
rect 37342 0 37454 800
rect 37986 0 38098 800
rect 39274 0 39386 800
rect 40562 0 40674 800
rect 41850 0 41962 800
rect 43138 0 43250 800
rect 44426 0 44538 800
rect 45714 0 45826 800
rect 47002 0 47114 800
rect 48290 0 48402 800
rect 49578 0 49690 800
rect 50866 0 50978 800
rect 52154 0 52266 800
rect 53442 0 53554 800
rect 54730 0 54842 800
rect 56018 0 56130 800
rect 56662 0 56774 800
rect 57950 0 58062 800
rect 59238 0 59350 800
rect 60526 0 60638 800
rect 61814 0 61926 800
rect 63102 0 63214 800
rect 64390 0 64502 800
rect 65678 0 65790 800
<< obsm2 >>
rect 802 67887 1866 68105
rect 2090 67887 3154 68105
rect 3378 67887 4442 68105
rect 4666 67887 5730 68105
rect 5954 67887 7018 68105
rect 7242 67887 8306 68105
rect 8530 67887 9594 68105
rect 9818 67887 10238 68105
rect 10462 67887 11526 68105
rect 11750 67887 12814 68105
rect 13038 67887 14102 68105
rect 14326 67887 15390 68105
rect 15614 67887 16678 68105
rect 16902 67887 17966 68105
rect 18190 67887 19254 68105
rect 19478 67887 20542 68105
rect 20766 67887 21830 68105
rect 22054 67887 23118 68105
rect 23342 67887 24406 68105
rect 24630 67887 25694 68105
rect 25918 67887 26982 68105
rect 27206 67887 28270 68105
rect 28494 67887 28914 68105
rect 29138 67887 30202 68105
rect 30426 67887 31490 68105
rect 31714 67887 32778 68105
rect 33002 67887 34066 68105
rect 34290 67887 35354 68105
rect 35578 67887 36642 68105
rect 36866 67887 37930 68105
rect 38154 67887 39218 68105
rect 39442 67887 40506 68105
rect 40730 67887 41794 68105
rect 42018 67887 43082 68105
rect 43306 67887 44370 68105
rect 44594 67887 45658 68105
rect 45882 67887 46946 68105
rect 47170 67887 47590 68105
rect 47814 67887 48878 68105
rect 49102 67887 50166 68105
rect 50390 67887 51454 68105
rect 51678 67887 52742 68105
rect 52966 67887 54030 68105
rect 54254 67887 55318 68105
rect 55542 67887 56606 68105
rect 56830 67887 57894 68105
rect 58118 67887 59182 68105
rect 59406 67887 60470 68105
rect 60694 67887 61758 68105
rect 61982 67887 63046 68105
rect 63270 67887 64334 68105
rect 64558 67887 65622 68105
rect 664 856 65760 67887
rect 802 734 1866 856
rect 2090 734 3154 856
rect 3378 734 4442 856
rect 4666 734 5730 856
rect 5954 734 7018 856
rect 7242 734 8306 856
rect 8530 734 9594 856
rect 9818 734 10882 856
rect 11106 734 12170 856
rect 12394 734 13458 856
rect 13682 734 14746 856
rect 14970 734 16034 856
rect 16258 734 17322 856
rect 17546 734 18610 856
rect 18834 734 19254 856
rect 19478 734 20542 856
rect 20766 734 21830 856
rect 22054 734 23118 856
rect 23342 734 24406 856
rect 24630 734 25694 856
rect 25918 734 26982 856
rect 27206 734 28270 856
rect 28494 734 29558 856
rect 29782 734 30846 856
rect 31070 734 32134 856
rect 32358 734 33422 856
rect 33646 734 34710 856
rect 34934 734 35998 856
rect 36222 734 37286 856
rect 37510 734 37930 856
rect 38154 734 39218 856
rect 39442 734 40506 856
rect 40730 734 41794 856
rect 42018 734 43082 856
rect 43306 734 44370 856
rect 44594 734 45658 856
rect 45882 734 46946 856
rect 47170 734 48234 856
rect 48458 734 49522 856
rect 49746 734 50810 856
rect 51034 734 52098 856
rect 52322 734 53386 856
rect 53610 734 54674 856
rect 54898 734 55962 856
rect 56186 734 56606 856
rect 56830 734 57894 856
rect 58118 734 59182 856
rect 59406 734 60470 856
rect 60694 734 61758 856
rect 61982 734 63046 856
rect 63270 734 64334 856
rect 64558 734 65622 856
<< metal3 >>
rect 0 67948 800 68188
rect 65799 67268 66599 67508
rect 0 66588 800 66828
rect 65799 65908 66599 66148
rect 0 65228 800 65468
rect 65799 64548 66599 64788
rect 0 63868 800 64108
rect 65799 63188 66599 63428
rect 0 62508 800 62748
rect 65799 61828 66599 62068
rect 0 61148 800 61388
rect 65799 60468 66599 60708
rect 0 59788 800 60028
rect 0 59108 800 59348
rect 65799 59108 66599 59348
rect 0 57748 800 57988
rect 65799 57748 66599 57988
rect 0 56388 800 56628
rect 65799 56388 66599 56628
rect 0 55028 800 55268
rect 65799 55028 66599 55268
rect 0 53668 800 53908
rect 65799 53668 66599 53908
rect 0 52308 800 52548
rect 65799 52308 66599 52548
rect 0 50948 800 51188
rect 65799 50948 66599 51188
rect 0 49588 800 49828
rect 65799 49588 66599 49828
rect 0 48228 800 48468
rect 65799 48228 66599 48468
rect 65799 47548 66599 47788
rect 0 46868 800 47108
rect 65799 46188 66599 46428
rect 0 45508 800 45748
rect 65799 44828 66599 45068
rect 0 44148 800 44388
rect 65799 43468 66599 43708
rect 0 42788 800 43028
rect 65799 42108 66599 42348
rect 0 41428 800 41668
rect 65799 40748 66599 40988
rect 0 40068 800 40308
rect 0 39388 800 39628
rect 65799 39388 66599 39628
rect 0 38028 800 38268
rect 65799 38028 66599 38268
rect 0 36668 800 36908
rect 65799 36668 66599 36908
rect 0 35308 800 35548
rect 65799 35308 66599 35548
rect 0 33948 800 34188
rect 65799 33948 66599 34188
rect 0 32588 800 32828
rect 65799 32588 66599 32828
rect 0 31228 800 31468
rect 65799 31228 66599 31468
rect 0 29868 800 30108
rect 65799 29868 66599 30108
rect 0 28508 800 28748
rect 65799 28508 66599 28748
rect 65799 27828 66599 28068
rect 0 27148 800 27388
rect 65799 26468 66599 26708
rect 0 25788 800 26028
rect 65799 25108 66599 25348
rect 0 24428 800 24668
rect 65799 23748 66599 23988
rect 0 23068 800 23308
rect 65799 22388 66599 22628
rect 0 21708 800 21948
rect 65799 21028 66599 21268
rect 0 20348 800 20588
rect 0 19668 800 19908
rect 65799 19668 66599 19908
rect 0 18308 800 18548
rect 65799 18308 66599 18548
rect 0 16948 800 17188
rect 65799 16948 66599 17188
rect 0 15588 800 15828
rect 65799 15588 66599 15828
rect 0 14228 800 14468
rect 65799 14228 66599 14468
rect 0 12868 800 13108
rect 65799 12868 66599 13108
rect 0 11508 800 11748
rect 65799 11508 66599 11748
rect 0 10148 800 10388
rect 65799 10148 66599 10388
rect 0 8788 800 9028
rect 65799 8788 66599 9028
rect 65799 8108 66599 8348
rect 0 7428 800 7668
rect 65799 6748 66599 6988
rect 0 6068 800 6308
rect 65799 5388 66599 5628
rect 0 4708 800 4948
rect 65799 4028 66599 4268
rect 0 3348 800 3588
rect 65799 2668 66599 2908
rect 0 1988 800 2228
rect 65799 1308 66599 1548
rect 0 628 800 868
rect 65799 -52 66599 188
<< obsm3 >>
rect 880 67868 65799 68101
rect 800 67588 65799 67868
rect 800 67188 65719 67588
rect 800 66908 65799 67188
rect 880 66508 65799 66908
rect 800 66228 65799 66508
rect 800 65828 65719 66228
rect 800 65548 65799 65828
rect 880 65148 65799 65548
rect 800 64868 65799 65148
rect 800 64468 65719 64868
rect 800 64188 65799 64468
rect 880 63788 65799 64188
rect 800 63508 65799 63788
rect 800 63108 65719 63508
rect 800 62828 65799 63108
rect 880 62428 65799 62828
rect 800 62148 65799 62428
rect 800 61748 65719 62148
rect 800 61468 65799 61748
rect 880 61068 65799 61468
rect 800 60788 65799 61068
rect 800 60388 65719 60788
rect 800 60108 65799 60388
rect 880 59708 65799 60108
rect 800 59428 65799 59708
rect 880 59028 65719 59428
rect 800 58068 65799 59028
rect 880 57668 65719 58068
rect 800 56708 65799 57668
rect 880 56308 65719 56708
rect 800 55348 65799 56308
rect 880 54948 65719 55348
rect 800 53988 65799 54948
rect 880 53588 65719 53988
rect 800 52628 65799 53588
rect 880 52228 65719 52628
rect 800 51268 65799 52228
rect 880 50868 65719 51268
rect 800 49908 65799 50868
rect 880 49508 65719 49908
rect 800 48548 65799 49508
rect 880 48148 65719 48548
rect 800 47868 65799 48148
rect 800 47468 65719 47868
rect 800 47188 65799 47468
rect 880 46788 65799 47188
rect 800 46508 65799 46788
rect 800 46108 65719 46508
rect 800 45828 65799 46108
rect 880 45428 65799 45828
rect 800 45148 65799 45428
rect 800 44748 65719 45148
rect 800 44468 65799 44748
rect 880 44068 65799 44468
rect 800 43788 65799 44068
rect 800 43388 65719 43788
rect 800 43108 65799 43388
rect 880 42708 65799 43108
rect 800 42428 65799 42708
rect 800 42028 65719 42428
rect 800 41748 65799 42028
rect 880 41348 65799 41748
rect 800 41068 65799 41348
rect 800 40668 65719 41068
rect 800 40388 65799 40668
rect 880 39988 65799 40388
rect 800 39708 65799 39988
rect 880 39308 65719 39708
rect 800 38348 65799 39308
rect 880 37948 65719 38348
rect 800 36988 65799 37948
rect 880 36588 65719 36988
rect 800 35628 65799 36588
rect 880 35228 65719 35628
rect 800 34268 65799 35228
rect 880 33868 65719 34268
rect 800 32908 65799 33868
rect 880 32508 65719 32908
rect 800 31548 65799 32508
rect 880 31148 65719 31548
rect 800 30188 65799 31148
rect 880 29788 65719 30188
rect 800 28828 65799 29788
rect 880 28428 65719 28828
rect 800 28148 65799 28428
rect 800 27748 65719 28148
rect 800 27468 65799 27748
rect 880 27068 65799 27468
rect 800 26788 65799 27068
rect 800 26388 65719 26788
rect 800 26108 65799 26388
rect 880 25708 65799 26108
rect 800 25428 65799 25708
rect 800 25028 65719 25428
rect 800 24748 65799 25028
rect 880 24348 65799 24748
rect 800 24068 65799 24348
rect 800 23668 65719 24068
rect 800 23388 65799 23668
rect 880 22988 65799 23388
rect 800 22708 65799 22988
rect 800 22308 65719 22708
rect 800 22028 65799 22308
rect 880 21628 65799 22028
rect 800 21348 65799 21628
rect 800 20948 65719 21348
rect 800 20668 65799 20948
rect 880 20268 65799 20668
rect 800 19988 65799 20268
rect 880 19588 65719 19988
rect 800 18628 65799 19588
rect 880 18228 65719 18628
rect 800 17268 65799 18228
rect 880 16868 65719 17268
rect 800 15908 65799 16868
rect 880 15508 65719 15908
rect 800 14548 65799 15508
rect 880 14148 65719 14548
rect 800 13188 65799 14148
rect 880 12788 65719 13188
rect 800 11828 65799 12788
rect 880 11428 65719 11828
rect 800 10468 65799 11428
rect 880 10068 65719 10468
rect 800 9108 65799 10068
rect 880 8708 65719 9108
rect 800 8428 65799 8708
rect 800 8028 65719 8428
rect 800 7748 65799 8028
rect 880 7348 65799 7748
rect 800 7068 65799 7348
rect 800 6668 65719 7068
rect 800 6388 65799 6668
rect 880 5988 65799 6388
rect 800 5708 65799 5988
rect 800 5308 65719 5708
rect 800 5028 65799 5308
rect 880 4628 65799 5028
rect 800 4348 65799 4628
rect 800 3948 65719 4348
rect 800 3668 65799 3948
rect 880 3268 65799 3668
rect 800 2988 65799 3268
rect 800 2588 65719 2988
rect 800 2308 65799 2588
rect 880 1908 65799 2308
rect 800 1628 65799 1908
rect 800 1395 65719 1628
<< metal4 >>
rect 4208 2128 4528 66416
rect 19568 2128 19888 66416
rect 34928 2128 35248 66416
rect 50288 2128 50608 66416
<< obsm4 >>
rect 10179 24787 19488 59397
rect 19968 24787 34717 59397
<< labels >>
rlabel metal3 s 0 62508 800 62748 6 active
port 1 nsew signal input
rlabel metal2 s 20598 0 20710 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 36698 67943 36810 68743 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 0 67948 800 68188 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 65799 57748 66599 57988 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 32190 0 32302 800 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 24462 67943 24574 68743 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 65799 60468 66599 60708 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 65799 6748 66599 6988 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 12870 67943 12982 68743 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 15446 67943 15558 68743 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 57950 0 58062 800 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 0 21708 800 21948 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 0 39388 800 39628 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 65799 22388 66599 22628 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 11582 67943 11694 68743 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 8362 67943 8474 68743 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 50866 0 50978 800 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 49578 0 49690 800 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 65799 15588 66599 15828 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 44426 0 44538 800 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 66322 67943 66434 68743 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 65799 27828 66599 28068 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 59788 800 60028 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 41850 0 41962 800 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 50222 67943 50334 68743 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 57950 67943 58062 68743 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 65799 43468 66599 43708 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 59238 67943 59350 68743 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 37986 67943 38098 68743 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 65799 42108 66599 42348 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 65799 65908 66599 66148 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 41428 800 41668 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 65799 46188 66599 46428 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 10294 67943 10406 68743 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 36054 0 36166 800 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 23068 800 23308 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 65799 39388 66599 39628 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 65799 21028 66599 21268 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 65799 19668 66599 19908 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 6068 800 6308 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 18022 67943 18134 68743 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 65799 4028 66599 4268 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 18666 0 18778 800 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 47646 67943 47758 68743 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 19310 67943 19422 68743 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 53442 0 53554 800 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 65799 29868 66599 30108 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 1922 67943 2034 68743 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 7074 0 7186 800 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 32834 67943 32946 68743 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 34122 67943 34234 68743 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 64390 0 64502 800 6 io_oeb[25]
port 57 nsew signal output
rlabel metal3 s 65799 53668 66599 53908 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 39274 67943 39386 68743 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 56662 0 56774 800 6 io_oeb[28]
port 60 nsew signal output
rlabel metal3 s 65799 44828 66599 45068 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 55374 67943 55486 68743 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 3210 67943 3322 68743 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 56018 0 56130 800 6 io_oeb[31]
port 64 nsew signal output
rlabel metal3 s 0 33948 800 34188 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 65678 0 65790 800 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 14158 67943 14270 68743 6 io_oeb[34]
port 67 nsew signal output
rlabel metal3 s 0 29868 800 30108 6 io_oeb[35]
port 68 nsew signal output
rlabel metal3 s 0 15588 800 15828 6 io_oeb[36]
port 69 nsew signal output
rlabel metal3 s 0 24428 800 24668 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 34766 0 34878 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 65799 1308 66599 1548 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 44148 800 44388 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 65799 25108 66599 25348 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 16734 67943 16846 68743 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 5786 0 5898 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 14802 0 14914 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 65799 64548 66599 64788 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 65799 38028 66599 38268 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 0 3348 800 3588 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 0 10148 800 10388 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 54730 0 54842 800 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 65799 55028 66599 55268 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 0 56388 800 56628 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 65799 36668 66599 36908 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 61814 67943 61926 68743 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 63102 0 63214 800 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 0 32588 800 32828 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 44426 67943 44538 68743 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 54086 67943 54198 68743 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 0 55028 800 55268 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 43138 0 43250 800 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 65799 31228 66599 31468 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 37342 0 37454 800 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 48934 67943 49046 68743 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 0 7428 800 7668 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 51510 67943 51622 68743 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 23174 0 23286 800 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 65799 2668 66599 2908 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 9650 0 9762 800 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 0 8788 800 9028 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 0 19668 800 19908 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 0 63868 800 64108 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 65799 10148 66599 10388 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 65799 56388 66599 56628 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 65799 52308 66599 52548 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 20598 67943 20710 68743 6 io_out[36]
port 107 nsew signal output
rlabel metal3 s 65799 61828 66599 62068 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 0 59108 800 59348 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 65799 40748 66599 40988 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 30258 67943 30370 68743 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 64390 67943 64502 68743 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 0 27148 800 27388 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 25750 0 25862 800 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 0 20348 800 20588 6 io_out[9]
port 115 nsew signal output
rlabel metal3 s 65799 11508 66599 11748 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal3 s 65799 8788 66599 9028 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal3 s 0 50948 800 51188 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 45714 0 45826 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal3 s 0 18308 800 18548 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 21886 67943 21998 68743 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 41850 67943 41962 68743 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 31546 67943 31658 68743 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 59238 0 59350 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 23174 67943 23286 68743 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal3 s 0 49588 800 49828 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 65678 67943 65790 68743 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal3 s 65799 12868 66599 13108 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal3 s 0 52308 800 52548 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 65799 5388 66599 5628 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 634 67943 746 68743 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 52154 0 52266 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal3 s 0 42788 800 43028 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 56662 67943 56774 68743 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal3 s 65799 33948 66599 34188 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 25750 67943 25862 68743 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 27038 67943 27150 68743 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal3 s 0 46868 800 47108 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal3 s 65799 16948 66599 17188 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 30902 0 31014 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal3 s 65799 63188 66599 63428 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 5786 67943 5898 68743 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 35410 67943 35522 68743 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal3 s 0 1988 800 2228 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal3 s 65799 23748 66599 23988 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal3 s 65799 49588 66599 49828 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 7074 67943 7186 68743 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal3 s 65799 35308 66599 35548 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal3 s 0 61148 800 61388 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal3 s 0 14228 800 14468 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal3 s 65799 59108 66599 59348 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 40562 67943 40674 68743 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 17378 0 17490 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal3 s 65799 26468 66599 26708 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal3 s 0 4708 800 4948 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal3 s 65799 8108 66599 8348 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal3 s 0 65228 800 65468 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 60526 0 60638 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 8362 0 8474 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 28326 0 28438 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal3 s 65799 18308 66599 18548 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal3 s 65799 67268 66599 67508 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal3 s 0 12868 800 13108 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 61814 0 61926 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 4498 0 4610 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal3 s 65799 28508 66599 28748 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal3 s 65799 50948 66599 51188 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 63102 67943 63214 68743 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 65799 -52 66599 188 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal2 s 60526 67943 60638 68743 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal2 s 40562 0 40674 800 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 48290 0 48402 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal2 s 4498 67943 4610 68743 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 28970 67943 29082 68743 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 36668 800 36908 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal2 s 12226 0 12338 800 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 3210 0 3322 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 43138 67943 43250 68743 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 28326 67943 28438 68743 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 52798 67943 52910 68743 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 65799 14228 66599 14468 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 0 53668 800 53908 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 65799 48228 66599 48468 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal2 s 13514 0 13626 800 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 24462 0 24574 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 65799 47548 66599 47788 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal2 s 37986 0 38098 800 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 47002 67943 47114 68743 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 45714 67943 45826 68743 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 66588 800 66828 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal2 s 9650 67943 9762 68743 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 47002 0 47114 800 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 57748 800 57988 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 66416 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 66416 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 66416 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 2128 50608 66416 6 vssd1
port 213 nsew ground input
rlabel metal3 s 65799 32588 66599 32828 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 66599 68743
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9347676
string GDS_FILE /home/proppy/src/github.com/mattvenn/wrapped_rgb_mixer/runs/RUN_2022.03.19_15.21.20/results/finishing/wrapped_rgb_mixer.magic.gds
string GDS_START 1237104
<< end >>

