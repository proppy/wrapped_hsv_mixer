* NGSPICE file created from wrapped_hsv_mixer.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt wrapped_hsv_mixer active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6524__106 vssd1 vssd1 vccd1 vccd1 _6524__106/HI _6632_/A sky130_fd_sc_hd__conb_1
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _5290_/A vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__buf_2
XFILLER_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5727_ _5727_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5727_/Y sky130_fd_sc_hd__nand2_1
X_5658_ _5731_/A _5731_/B _5657_/Y vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__o21a_1
X_5589_ _5647_/A _5622_/A _5622_/B _5588_/X vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__o31ai_4
X_4609_ _4525_/A _4523_/X _4530_/X _4531_/Y _4608_/X vssd1 vssd1 vccd1 vccd1 _4609_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4960_ _4960_/A _4960_/B vssd1 vssd1 vccd1 vccd1 _5231_/C sky130_fd_sc_hd__nor2_1
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3911_ _5287_/A vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__clkbuf_2
X_4891_ _4891_/A _4891_/B _4891_/C _4891_/D vssd1 vssd1 vccd1 vccd1 _4899_/A sky130_fd_sc_hd__nand4_1
X_3842_ _3843_/A _3843_/B _3843_/C vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__o21ai_1
X_6630_ _6630_/A _3329_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_6561_ _6561_/A _3247_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3773_ _3483_/A _3518_/A _3482_/X vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__o21ba_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _6318_/Q _5487_/B _5471_/B _5487_/A vssd1 vssd1 vccd1 vccd1 _5512_/X sky130_fd_sc_hd__a22o_1
X_5443_ _5443_/A _5443_/B vssd1 vssd1 vccd1 vccd1 _5470_/B sky130_fd_sc_hd__nor2_2
X_5374_ _5411_/A _5411_/B _5373_/X vssd1 vssd1 vccd1 vccd1 _5376_/B sky130_fd_sc_hd__o21ai_2
X_4325_ _4461_/B _4325_/B vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__xnor2_4
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4391_/B _4391_/C vssd1 vssd1 vccd1 vccd1 _4256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4187_ _4387_/B vssd1 vssd1 vccd1 vccd1 _4424_/B sky130_fd_sc_hd__buf_2
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6517__99 vssd1 vssd1 vccd1 vccd1 _6517__99/HI _6625_/A sky130_fd_sc_hd__conb_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4110_ _4110_/A _4110_/B _4144_/A vssd1 vssd1 vccd1 vccd1 _4148_/B sky130_fd_sc_hd__or3_1
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5090_ _5090_/A _5090_/B _5090_/C vssd1 vssd1 vccd1 vccd1 _5091_/B sky130_fd_sc_hd__nor3_1
X_4041_ _5712_/A _4041_/B _4047_/A _4041_/D vssd1 vssd1 vccd1 vccd1 _4047_/B sky130_fd_sc_hd__nand4_1
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5992_ _6010_/B vssd1 vssd1 vccd1 vccd1 _5992_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4943_ _4623_/A _4924_/B _4929_/B _4928_/A vssd1 vssd1 vccd1 vccd1 _4943_/X sky130_fd_sc_hd__a31o_1
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4874_ _4874_/A _4886_/B _4874_/C vssd1 vssd1 vccd1 vccd1 _4875_/B sky130_fd_sc_hd__and3_1
XFILLER_60_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6613_ _6613_/A _3305_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_3825_ _4383_/A vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__clkbuf_2
X_6544_ _6544_/A _3227_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_3756_ _4131_/A _4185_/A vssd1 vssd1 vccd1 vccd1 _4101_/C sky130_fd_sc_hd__nor2_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5426_ _5386_/A _5455_/B _5455_/C _5458_/B _5387_/A vssd1 vssd1 vccd1 vccd1 _5426_/X
+ sky130_fd_sc_hd__a32o_1
X_3687_ _3690_/A _3690_/C _3706_/A vssd1 vssd1 vccd1 vccd1 _3692_/A sky130_fd_sc_hd__o21ai_1
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5357_ _5359_/A _5359_/B _5355_/A vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__o21ai_4
XFILLER_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5288_ _5288_/A _5288_/B vssd1 vssd1 vccd1 vccd1 _5289_/B sky130_fd_sc_hd__nand2_1
X_4308_ _4308_/A _4308_/B vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__xnor2_1
X_4239_ _4265_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4239_/X sky130_fd_sc_hd__or2_1
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _4557_/A _4557_/B _4565_/X _4589_/X vssd1 vssd1 vccd1 vccd1 _4590_/X sky130_fd_sc_hd__a22o_1
X_3610_ _4755_/B _3566_/A _3570_/C _4659_/B vssd1 vssd1 vccd1 vccd1 _3610_/X sky130_fd_sc_hd__a22o_1
X_3541_ _3591_/A _3591_/B vssd1 vssd1 vccd1 vccd1 _3547_/B sky130_fd_sc_hd__nand2_1
X_3472_ _6342_/Q _3472_/B vssd1 vssd1 vccd1 vccd1 _3473_/B sky130_fd_sc_hd__nor2_1
X_6260_ _6280_/A _6260_/B vssd1 vssd1 vccd1 vccd1 _6260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5211_ _5211_/A _5240_/B vssd1 vssd1 vccd1 vccd1 _5222_/A sky130_fd_sc_hd__nand2_1
X_6191_ _6191_/A vssd1 vssd1 vccd1 vccd1 _6379_/D sky130_fd_sc_hd__clkbuf_1
X_5142_ _5142_/A _5141_/A vssd1 vssd1 vccd1 vccd1 _5142_/X sky130_fd_sc_hd__or2b_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5073_ _5134_/A _5134_/B _5072_/Y vssd1 vssd1 vccd1 vccd1 _5081_/B sky130_fd_sc_hd__o21ai_2
X_4024_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _4025_/C sky130_fd_sc_hd__xor2_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5975_ _5981_/A _6014_/A _5911_/X vssd1 vssd1 vccd1 vccd1 _5975_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4926_ _4927_/A _4927_/B vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__and2_1
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4857_ _4863_/A _4857_/B vssd1 vssd1 vccd1 vccd1 _4858_/C sky130_fd_sc_hd__xnor2_1
X_3808_ _3808_/A _3808_/B vssd1 vssd1 vccd1 vccd1 _3822_/B sky130_fd_sc_hd__xor2_1
X_4788_ _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4794_/C sky130_fd_sc_hd__nor2_1
X_3739_ _4814_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _4957_/C sky130_fd_sc_hd__nand2_2
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _5373_/B _5406_/Y _5408_/X vssd1 vssd1 vccd1 vccd1 _5440_/B sky130_fd_sc_hd__o21ai_2
X_6389_ _6396_/CLK _6389_/D vssd1 vssd1 vccd1 vccd1 _6389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6501__83 vssd1 vssd1 vccd1 vccd1 _6501__83/HI _6609_/A sky130_fd_sc_hd__conb_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5760_ _5823_/B _5758_/Y _5868_/B _5759_/Y vssd1 vssd1 vccd1 vccd1 _5760_/X sky130_fd_sc_hd__a22o_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4711_/A _4711_/B _4872_/B _4711_/D vssd1 vssd1 vccd1 vccd1 _4713_/A sky130_fd_sc_hd__and4_1
X_5691_ _5691_/A _5691_/B vssd1 vssd1 vccd1 vccd1 _5691_/Y sky130_fd_sc_hd__xnor2_1
X_4642_ _6340_/Q _4660_/B _4648_/B _4642_/D vssd1 vssd1 vccd1 vccd1 _4751_/C sky130_fd_sc_hd__or4_4
X_4573_ _4573_/A _4573_/B vssd1 vssd1 vccd1 vccd1 _5560_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3524_ _4697_/B _3522_/X _3523_/X vssd1 vssd1 vccd1 vccd1 _3546_/A sky130_fd_sc_hd__a21bo_1
X_6312_ _6425_/Q _6310_/B _6007_/X vssd1 vssd1 vccd1 vccd1 _6312_/Y sky130_fd_sc_hd__a21oi_1
X_6243_ _6399_/Q _6243_/B vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__and2_1
X_3455_ _4660_/B vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3386_ _6332_/Q vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__clkbuf_2
X_6174_ _6174_/A vssd1 vssd1 vccd1 vccd1 _6373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5125_ _5125_/A _5125_/B vssd1 vssd1 vccd1 vccd1 _5126_/B sky130_fd_sc_hd__xnor2_2
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5056_ _5092_/A _5092_/B vssd1 vssd1 vccd1 vccd1 _5057_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4007_ _3978_/A _3978_/B _3978_/C vssd1 vssd1 vccd1 vccd1 _4027_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5958_ input8/X vssd1 vssd1 vccd1 vccd1 _6282_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4909_ _4909_/A _4909_/B _4909_/C vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5889_ _6422_/Q _5885_/X _5888_/Y _6423_/Q vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3241_/A vssd1 vssd1 vccd1 vccd1 _3240_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5812_ input8/X vssd1 vssd1 vccd1 vccd1 _6310_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5743_ _5743_/A vssd1 vssd1 vccd1 vccd1 _5743_/X sky130_fd_sc_hd__clkbuf_2
X_5674_ _5674_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__xnor2_1
X_4625_ _4688_/B vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__clkbuf_4
X_4556_ _5937_/A _4558_/B _4555_/X vssd1 vssd1 vccd1 vccd1 _4557_/B sky130_fd_sc_hd__a21o_1
X_3507_ _3507_/A _3507_/B vssd1 vssd1 vccd1 vccd1 _3515_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4487_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _5789_/A sky130_fd_sc_hd__xor2_4
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3438_ _3438_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3446_/C sky130_fd_sc_hd__xnor2_1
XFILLER_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6226_ _6224_/X _6225_/X _6334_/D vssd1 vssd1 vccd1 vccd1 _6226_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3369_ _5159_/A vssd1 vssd1 vccd1 vccd1 _5102_/A sky130_fd_sc_hd__clkbuf_2
X_6157_ _6100_/X _6152_/X _6153_/X _6156_/X vssd1 vssd1 vccd1 vccd1 _6365_/D sky130_fd_sc_hd__a31o_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5282_/A _5288_/B vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__nand2_2
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6492__74 vssd1 vssd1 vccd1 vccd1 _6492__74/HI _6600_/A sky130_fd_sc_hd__conb_1
X_6088_ _6104_/B _6088_/B vssd1 vssd1 vccd1 vccd1 _6089_/B sky130_fd_sc_hd__or2_1
X_5039_ _5039_/A _5039_/B vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4410_ _5560_/A _4412_/B _4413_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__a31o_1
X_5390_ _5390_/A _5390_/B vssd1 vssd1 vccd1 vccd1 _5390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4341_ _4341_/A _4341_/B vssd1 vssd1 vccd1 vccd1 _4347_/C sky130_fd_sc_hd__xnor2_4
X_4272_ _4272_/A _4272_/B _4336_/A vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__and3_1
X_3223_ input1/X vssd1 vssd1 vccd1 vccd1 _3248_/A sky130_fd_sc_hd__buf_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6011_ _4630_/C _6010_/B _6004_/X vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ _5324_/A vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5726_ _5726_/A _5726_/B vssd1 vssd1 vccd1 vccd1 _5729_/B sky130_fd_sc_hd__xnor2_1
X_5657_ _5758_/A _5702_/A vssd1 vssd1 vccd1 vccd1 _5657_/Y sky130_fd_sc_hd__nand2_1
X_5588_ _5648_/A _5228_/A _5647_/A vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__a21o_1
X_4608_ _4606_/X _4607_/X _4528_/X _4529_/Y vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4539_ _4540_/A _4540_/B vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6209_ _6385_/Q _6213_/B vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__and2_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3910_ _5350_/A vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4890_ _3685_/A _4873_/B _4895_/D _4895_/A vssd1 vssd1 vccd1 vccd1 _4899_/B sky130_fd_sc_hd__a22o_1
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3841_ _3841_/A _3841_/B vssd1 vssd1 vccd1 vccd1 _3843_/C sky130_fd_sc_hd__xor2_1
X_3772_ _3804_/B _3805_/B _3771_/Y vssd1 vssd1 vccd1 vccd1 _3788_/B sky130_fd_sc_hd__a21o_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6560_ _6560_/A _3246_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
X_5511_ _5511_/A _5532_/A vssd1 vssd1 vccd1 vccd1 _5511_/Y sky130_fd_sc_hd__nor2_2
X_5442_ _6321_/Q _5471_/B _4272_/B vssd1 vssd1 vccd1 vccd1 _5443_/B sky130_fd_sc_hd__a21oi_1
X_5373_ _5373_/A _5373_/B vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__or2_1
X_4324_ _4326_/A _4326_/B _4323_/X vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__a21oi_2
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4255_ _4255_/A vssd1 vssd1 vccd1 vccd1 _4391_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4186_ _4330_/B vssd1 vssd1 vccd1 vccd1 _4387_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6462__44 vssd1 vssd1 vccd1 vccd1 _6462__44/HI _6567_/A sky130_fd_sc_hd__conb_1
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5709_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5710_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4040_ _5121_/A _4079_/B _4022_/B _4037_/Y vssd1 vssd1 vccd1 vccd1 _4041_/D sky130_fd_sc_hd__a211o_1
XFILLER_77_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5991_ _5985_/A _5978_/A _5981_/A _6010_/B vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__a31o_1
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _4981_/S _4980_/A vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4873_ _4891_/A _4873_/B vssd1 vssd1 vccd1 vccd1 _4875_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6612_ _6612_/A _3307_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3824_ _6320_/Q vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__clkbuf_2
X_3755_ _4184_/A _4184_/B vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__and2_1
X_6543_ _6543_/A _3226_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3686_ _3705_/B _3705_/C _3705_/A vssd1 vssd1 vccd1 vccd1 _3706_/A sky130_fd_sc_hd__a21o_1
X_5425_ _5425_/A _5492_/B _5492_/C vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__and3_1
X_5356_ _5356_/A _5514_/B vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__nand2_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5287_ _5287_/A _5392_/B vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__nand2_1
X_4307_ _4307_/A _4387_/B vssd1 vssd1 vccd1 vccd1 _4308_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4238_ _4238_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4169_ _4212_/A _5322_/A _4169_/C _4340_/B vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__and4_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3540_ _4800_/A _3685_/B vssd1 vssd1 vccd1 vccd1 _3591_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5210_ _5210_/A _5210_/B vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__xnor2_2
X_3471_ _6331_/Q vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__inv_2
X_6190_ _6378_/Q _6194_/B vssd1 vssd1 vccd1 vccd1 _6191_/A sky130_fd_sc_hd__and2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5141_ _5141_/A _5142_/A vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__xnor2_1
X_5072_ _5072_/A _5072_/B vssd1 vssd1 vccd1 vccd1 _5072_/Y sky130_fd_sc_hd__nand2_1
X_4023_ _4022_/A _4022_/B _3974_/A _3969_/X vssd1 vssd1 vccd1 vccd1 _4025_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6432__14 vssd1 vssd1 vccd1 vccd1 _6432__14/HI _6537_/A sky130_fd_sc_hd__conb_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5974_ _6014_/A vssd1 vssd1 vccd1 vccd1 _5982_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4925_ _3466_/A _4820_/B _4716_/X _4710_/A vssd1 vssd1 vccd1 vccd1 _4927_/B sky130_fd_sc_hd__a22o_1
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4856_ _4862_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4857_/B sky130_fd_sc_hd__xnor2_1
X_3807_ _5356_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__nand2_1
X_4787_ _4787_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__xnor2_1
X_3738_ _4895_/A vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3669_ _3669_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _3670_/B sky130_fd_sc_hd__xnor2_2
X_5408_ _5367_/A _5533_/B _5545_/B _5316_/A vssd1 vssd1 vccd1 vccd1 _5408_/X sky130_fd_sc_hd__a22o_1
X_6388_ _6388_/CLK _6388_/D vssd1 vssd1 vccd1 vccd1 _6388_/Q sky130_fd_sc_hd__dfxtp_1
X_5339_ _5331_/B _5339_/B vssd1 vssd1 vccd1 vccd1 _5339_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6498__80 vssd1 vssd1 vccd1 vccd1 _6498__80/HI _6606_/A sky130_fd_sc_hd__conb_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4710_ _4710_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__nand2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5723_/A _5723_/B vssd1 vssd1 vccd1 vccd1 _5690_/Y sky130_fd_sc_hd__nor2_1
X_4641_ _4660_/C vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__clkbuf_2
X_4572_ _4572_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4596_/C sky130_fd_sc_hd__xnor2_4
X_3523_ _4763_/A _3699_/C _3685_/B _4673_/B vssd1 vssd1 vccd1 vccd1 _3523_/X sky130_fd_sc_hd__a22o_1
X_6311_ _6424_/Q _6307_/B _6310_/Y vssd1 vssd1 vccd1 vccd1 _6424_/D sky130_fd_sc_hd__o21a_1
X_6242_ _6242_/A vssd1 vssd1 vccd1 vccd1 _6399_/D sky130_fd_sc_hd__clkbuf_1
X_3454_ _6346_/Q _6345_/Q _6339_/Q vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__a21o_2
X_3385_ _4630_/A _3395_/B vssd1 vssd1 vccd1 vccd1 _3385_/Y sky130_fd_sc_hd__nand2_1
X_6173_ _6372_/Q _6183_/B vssd1 vssd1 vccd1 vccd1 _6174_/A sky130_fd_sc_hd__and2_1
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _5124_/A _5124_/B vssd1 vssd1 vccd1 vccd1 _5125_/B sky130_fd_sc_hd__xnor2_4
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5055_ _5055_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5057_/A sky130_fd_sc_hd__nor2_2
X_4006_ _4005_/B _4005_/C _4005_/A vssd1 vssd1 vccd1 vccd1 _4474_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5957_ _5851_/X _5951_/X _5950_/B vssd1 vssd1 vccd1 vccd1 _5957_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4908_ _4955_/B _5275_/B _5275_/A vssd1 vssd1 vccd1 vccd1 _4953_/C sky130_fd_sc_hd__o21a_1
X_5888_ _5945_/A _5870_/X _5887_/X _5807_/X vssd1 vssd1 vccd1 vccd1 _5888_/Y sky130_fd_sc_hd__a22oi_2
X_4839_ _4839_/A _4861_/A vssd1 vssd1 vccd1 vccd1 _4841_/A sky130_fd_sc_hd__nand2_2
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5811_ _5802_/X _5809_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5742_ _5742_/A _5742_/B vssd1 vssd1 vccd1 vccd1 _5742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5673_ _5673_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5675_/B sky130_fd_sc_hd__xor2_2
X_4624_ _4624_/A vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ _4554_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__and2b_1
X_3506_ _3506_/A _3501_/B vssd1 vssd1 vccd1 vccd1 _3507_/B sky130_fd_sc_hd__or2b_1
X_4486_ _4486_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _5805_/A sky130_fd_sc_hd__xnor2_4
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3437_ _3438_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3440_/B sky130_fd_sc_hd__nor2_1
X_6225_ _6389_/Q _6388_/Q _6391_/Q _6390_/Q vssd1 vssd1 vccd1 vccd1 _6225_/X sky130_fd_sc_hd__or4_1
X_3368_ _4109_/A vssd1 vssd1 vccd1 vccd1 _5159_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6156_ _6358_/Q _6357_/Q _6155_/X _6325_/D vssd1 vssd1 vccd1 vccd1 _6156_/X sky130_fd_sc_hd__o31a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5107_ _5428_/B vssd1 vssd1 vccd1 vccd1 _5288_/B sky130_fd_sc_hd__buf_2
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3299_ _3303_/A vssd1 vssd1 vccd1 vccd1 _3299_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6087_ _6104_/B _6103_/B vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5038_ _5038_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5039_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6468__50 vssd1 vssd1 vccd1 vccd1 _6468__50/HI _6573_/A sky130_fd_sc_hd__conb_1
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _5425_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4341_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4271_ _5950_/A _4573_/B vssd1 vssd1 vccd1 vccd1 _4272_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3222_ _3222_/A vssd1 vssd1 vccd1 vccd1 _3222_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6010_ _6010_/A _6010_/B vssd1 vssd1 vccd1 vccd1 _6013_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3986_ _5362_/A vssd1 vssd1 vccd1 vccd1 _5324_/A sky130_fd_sc_hd__clkbuf_2
X_5725_ _5672_/Y _5676_/X _5677_/Y _5683_/X _5724_/X vssd1 vssd1 vccd1 vccd1 _5729_/A
+ sky130_fd_sc_hd__a221oi_1
X_5656_ _5758_/A _5702_/A vssd1 vssd1 vccd1 vccd1 _5731_/B sky130_fd_sc_hd__nor2_1
X_4607_ _4607_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__or2_1
X_5587_ _5191_/B _5191_/C _5191_/A vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__a21o_1
XFILLER_117_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4538_ _4538_/A _4545_/A vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__xnor2_2
X_4469_ _4515_/A _4515_/B _4467_/Y _4468_/X vssd1 vssd1 vccd1 vccd1 _4469_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_89_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6208_ _6208_/A vssd1 vssd1 vccd1 vccd1 _6385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6139_ _6358_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__and2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _5851_/A _3849_/B vssd1 vssd1 vccd1 vccd1 _3841_/B sky130_fd_sc_hd__nand2_1
X_3771_ _3518_/B _3561_/A _3518_/A vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5510_ _6318_/Q _5510_/B vssd1 vssd1 vccd1 vccd1 _5532_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5441_ _5441_/A _5510_/B _5441_/C vssd1 vssd1 vccd1 vccd1 _5443_/A sky130_fd_sc_hd__and3_1
X_5372_ _5373_/A _5373_/B vssd1 vssd1 vccd1 vccd1 _5411_/B sky130_fd_sc_hd__xnor2_1
X_4323_ _4322_/B _4323_/B vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__and2b_1
X_6530__112 vssd1 vssd1 vccd1 vccd1 _6530__112/HI _6638_/A sky130_fd_sc_hd__conb_1
XFILLER_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4254_ _4254_/A vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4185_ _4185_/A _4185_/B vssd1 vssd1 vccd1 vccd1 _4330_/B sky130_fd_sc_hd__or2_1
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3969_ _3973_/B vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__clkbuf_2
X_5708_ _5709_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__and2_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5639_ _5639_/A _5639_/B vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__xnor2_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6438__20 vssd1 vssd1 vccd1 vccd1 _6438__20/HI _6543_/A sky130_fd_sc_hd__conb_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5990_ _5997_/B vssd1 vssd1 vccd1 vccd1 _6010_/B sky130_fd_sc_hd__clkbuf_2
X_4941_ _4941_/A _4941_/B vssd1 vssd1 vccd1 vccd1 _4980_/A sky130_fd_sc_hd__nand2_1
X_4872_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__nand2_1
X_3823_ _3835_/B _3835_/A vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__and2b_1
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6611_ _6611_/A _3309_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
X_3754_ _3754_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _4184_/B sky130_fd_sc_hd__xnor2_1
X_6542_ _6542_/A _3225_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_3685_ _3685_/A _3685_/B vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__nand2_1
X_5424_ _5424_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__and2_1
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5355_ _5355_/A _5355_/B vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__nand2_2
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4306_ _4306_/A _4306_/B vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5286_ _5292_/A _5292_/B vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__xor2_2
X_4237_ _4237_/A _4237_/B vssd1 vssd1 vccd1 vccd1 _4265_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4212_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4168_/X sky130_fd_sc_hd__and2_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4099_ _5159_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3470_ _3477_/A _3470_/B vssd1 vssd1 vccd1 vccd1 _3484_/B sky130_fd_sc_hd__or2_1
XFILLER_108_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5140_ _5140_/A _5140_/B vssd1 vssd1 vccd1 vccd1 _5142_/A sky130_fd_sc_hd__xnor2_1
XFILLER_111_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5071_ _5079_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _5134_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4022_ _4022_/A _4022_/B _3974_/A _3969_/X vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__or4bb_1
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5973_ _6001_/S vssd1 vssd1 vccd1 vccd1 _6014_/A sky130_fd_sc_hd__clkbuf_2
X_4924_ _4924_/A _4924_/B vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _4855_/A _4855_/B _4855_/C vssd1 vssd1 vccd1 vccd1 _4856_/B sky130_fd_sc_hd__and3_1
X_3806_ _3973_/B vssd1 vssd1 vccd1 vccd1 _4154_/B sky130_fd_sc_hd__buf_2
X_4786_ _4786_/A vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__inv_2
X_3737_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__buf_2
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3668_ _3765_/B _3668_/B vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__xnor2_4
X_3599_ _3600_/B _3599_/B vssd1 vssd1 vccd1 vccd1 _3605_/B sky130_fd_sc_hd__xnor2_2
X_5407_ _5407_/A _5514_/B vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__nand2_1
X_6387_ _6388_/CLK _6387_/D vssd1 vssd1 vccd1 vccd1 _6387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5338_ _5338_/A _5338_/B vssd1 vssd1 vccd1 vccd1 _5358_/B sky130_fd_sc_hd__xnor2_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5269_ _5271_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _6346_/Q _6345_/Q _6338_/Q _6337_/Q _6336_/Q vssd1 vssd1 vccd1 vccd1 _4660_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_30_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6310_ _6310_/A _6310_/B vssd1 vssd1 vccd1 vccd1 _6310_/Y sky130_fd_sc_hd__nor2_1
X_4571_ _5697_/A _4571_/B vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__xor2_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3522_ _4763_/A _3699_/C _3685_/B vssd1 vssd1 vccd1 vccd1 _3522_/X sky130_fd_sc_hd__and3_1
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3453_ _3463_/A _3489_/A vssd1 vssd1 vccd1 vccd1 _3469_/B sky130_fd_sc_hd__or2_1
X_6241_ _6398_/Q _6243_/B vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__and2_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6172_ _6172_/A vssd1 vssd1 vccd1 vccd1 _6372_/D sky130_fd_sc_hd__clkbuf_1
X_5123_ _5004_/A _5004_/B _5095_/A vssd1 vssd1 vccd1 vccd1 _5124_/B sky130_fd_sc_hd__a21boi_2
XFILLER_97_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3384_ _3430_/B vssd1 vssd1 vccd1 vccd1 _3395_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5054_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__nor2_2
X_4005_ _4005_/A _4005_/B _4005_/C vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__nand3_1
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ _5851_/X _5842_/A _5951_/X _5950_/B vssd1 vssd1 vccd1 vccd1 _5956_/X sky130_fd_sc_hd__a31o_1
X_4907_ _4907_/A _4907_/B vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__xnor2_1
X_5887_ _5866_/X _5804_/X _5805_/X _5823_/C vssd1 vssd1 vccd1 vccd1 _5887_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4838_ _4839_/A _4838_/B _4838_/C vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4769_ _4956_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _4769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5810_ _6407_/Q _5808_/Y _5753_/X _6408_/Q vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5741_ _5803_/A _5748_/A _5803_/B _5634_/A vssd1 vssd1 vccd1 vccd1 _5742_/B sky130_fd_sc_hd__o31a_1
X_5672_ _5672_/A _5672_/B vssd1 vssd1 vccd1 vccd1 _5672_/Y sky130_fd_sc_hd__xnor2_1
X_4623_ _4623_/A vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4554_ _4554_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4558_/B sky130_fd_sc_hd__xnor2_1
XFILLER_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3505_ _3511_/A _3511_/B vssd1 vssd1 vccd1 vccd1 _3513_/A sky130_fd_sc_hd__or2b_1
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6224_ _6385_/Q _6384_/Q _6387_/Q _6386_/Q vssd1 vssd1 vccd1 vccd1 _6224_/X sky130_fd_sc_hd__or4_1
X_4485_ _4485_/A _3888_/X vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__or2b_2
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3436_ _3434_/A _3449_/A _3467_/A vssd1 vssd1 vccd1 vccd1 _3438_/B sky130_fd_sc_hd__o21a_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3367_ _5367_/A vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__clkbuf_2
X_6155_ _6360_/Q _6359_/Q _6155_/C vssd1 vssd1 vccd1 vccd1 _6155_/X sky130_fd_sc_hd__or3_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5106_/A _5106_/B vssd1 vssd1 vccd1 vccd1 _5428_/B sky130_fd_sc_hd__xnor2_4
X_6086_ _6343_/Q _6032_/X _6083_/X _6085_/Y _5948_/X vssd1 vssd1 vccd1 vccd1 _6343_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5037_ _5038_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__and2_1
X_3298_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3303_/A sky130_fd_sc_hd__buf_12
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5939_ _5785_/A _5933_/C _5931_/X vssd1 vssd1 vccd1 vccd1 _5940_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6483__65 vssd1 vssd1 vccd1 vccd1 _6483__65/HI _6591_/A sky130_fd_sc_hd__conb_1
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4270_ _4957_/B vssd1 vssd1 vccd1 vccd1 _4573_/B sky130_fd_sc_hd__buf_2
XFILLER_98_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3221_ _3222_/A vssd1 vssd1 vccd1 vccd1 _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3985_ _5425_/A vssd1 vssd1 vccd1 vccd1 _5362_/A sky130_fd_sc_hd__buf_2
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5724_ _5677_/Y _5683_/X _5690_/Y _5722_/X _5723_/Y vssd1 vssd1 vccd1 vccd1 _5724_/X
+ sky130_fd_sc_hd__o221a_1
X_5655_ _5655_/A _5655_/B vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__xor2_2
X_4606_ _4607_/A _4607_/B _4604_/A vssd1 vssd1 vccd1 vccd1 _4606_/X sky130_fd_sc_hd__a21bo_1
XFILLER_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5586_ _5617_/B _5619_/A _5619_/B _5585_/Y vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__a31oi_4
X_4537_ _4601_/A _4536_/C _5672_/A vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__a21o_1
X_4468_ _4205_/B _4468_/B vssd1 vssd1 vccd1 vccd1 _4468_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3419_ _4623_/A _3430_/C _3385_/Y vssd1 vssd1 vccd1 vccd1 _3441_/C sky130_fd_sc_hd__a21o_1
XFILLER_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6207_ _6384_/Q _6213_/B vssd1 vssd1 vccd1 vccd1 _6208_/A sky130_fd_sc_hd__and2_1
X_4399_ _4399_/A _4399_/B vssd1 vssd1 vccd1 vccd1 _4403_/B sky130_fd_sc_hd__xor2_4
X_6138_ _6138_/A vssd1 vssd1 vccd1 vccd1 _6358_/D sky130_fd_sc_hd__clkbuf_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6069_ _6077_/B _6068_/Y _6041_/A vssd1 vssd1 vccd1 vccd1 _6069_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3770_ _3813_/A _3813_/B _3564_/A vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__a21o_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5440_ _5440_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__xnor2_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5371_ _5371_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5373_/B sky130_fd_sc_hd__nand2_1
X_4322_ _4323_/B _4322_/B vssd1 vssd1 vccd1 vccd1 _4326_/B sky130_fd_sc_hd__xnor2_4
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4253_ _6320_/Q vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__inv_4
XFILLER_86_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4184_ _4184_/A _4184_/B vssd1 vssd1 vccd1 vccd1 _4185_/B sky130_fd_sc_hd__nor2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6425_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3968_ _5000_/A _4008_/B _4009_/B _3966_/Y vssd1 vssd1 vccd1 vccd1 _3977_/B sky130_fd_sc_hd__a31o_1
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5707_/A vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__inv_2
X_3899_ _5060_/A _3958_/B _4008_/B _5433_/A vssd1 vssd1 vccd1 vccd1 _3900_/B sky130_fd_sc_hd__a22oi_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5638_ _5654_/A _5654_/B _5596_/X vssd1 vssd1 vccd1 vccd1 _5639_/B sky130_fd_sc_hd__a21bo_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5569_ _5673_/A _5673_/B _5568_/Y vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6453__35 vssd1 vssd1 vccd1 vccd1 _6453__35/HI _6558_/A sky130_fd_sc_hd__conb_1
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _4936_/B _4937_/A _4977_/B _4939_/Y vssd1 vssd1 vccd1 vccd1 _4978_/B sky130_fd_sc_hd__o22a_1
X_4871_ _4871_/A _4871_/B vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__or2_1
X_3822_ _3822_/A _3822_/B vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6610_ _6610_/A _3312_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_20_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6541_ _6541_/A _3222_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _4814_/A _4904_/A _4957_/C _4802_/A vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__o22a_1
X_3684_ _3683_/A _3683_/B _3703_/B vssd1 vssd1 vccd1 vccd1 _3705_/C sky130_fd_sc_hd__a21o_1
X_5423_ _5545_/B vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__clkbuf_2
X_5354_ _5353_/A _5353_/B _5353_/C vssd1 vssd1 vccd1 vccd1 _5355_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _4305_/A _4305_/B vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5285_ _5237_/Y _5318_/A _5326_/A vssd1 vssd1 vccd1 vccd1 _5292_/B sky130_fd_sc_hd__o21ai_2
X_4236_ _4236_/A _4268_/A vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__nor2_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _4167_/A _4167_/B vssd1 vssd1 vccd1 vccd1 _4468_/B sky130_fd_sc_hd__and2_2
XFILLER_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4098_ _4114_/C _4098_/B vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5070_ _5137_/B _5070_/B vssd1 vssd1 vccd1 vccd1 _5071_/B sky130_fd_sc_hd__nand2_1
X_4021_ _5288_/A _4021_/B _4021_/C vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__and3_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5972_ _5968_/X _5969_/Y _5970_/X _5971_/X vssd1 vssd1 vccd1 vccd1 _6001_/S sky130_fd_sc_hd__o22a_2
X_4923_ _4732_/A _4923_/B vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__and2b_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4854_ _4891_/B _4854_/B vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__nand2_1
X_3805_ _3805_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__xor2_4
X_4785_ _5979_/A _4924_/B _4785_/C vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__and3_1
X_3736_ _3736_/A _3736_/B vssd1 vssd1 vccd1 vccd1 _3747_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3667_ _3670_/A _3665_/X _3666_/Y vssd1 vssd1 vccd1 vccd1 _3668_/B sky130_fd_sc_hd__a21boi_4
X_3598_ _3637_/A _3637_/B _3597_/X vssd1 vssd1 vccd1 vccd1 _3599_/B sky130_fd_sc_hd__o21ba_1
X_5406_ _5406_/A _5545_/B vssd1 vssd1 vccd1 vccd1 _5406_/Y sky130_fd_sc_hd__nand2_1
X_6386_ _6388_/CLK _6386_/D vssd1 vssd1 vccd1 vccd1 _6386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5337_ _5337_/A _5337_/B vssd1 vssd1 vccd1 vccd1 _5338_/B sky130_fd_sc_hd__or2_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _5268_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__xor2_2
XFILLER_85_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4219_ _5555_/C vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__buf_2
X_5199_ _5199_/A _5199_/B vssd1 vssd1 vccd1 vccd1 _5201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_18_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _5697_/A _4571_/B _4569_/Y vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__a21oi_1
X_3521_ _4886_/A vssd1 vssd1 vccd1 vccd1 _4688_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3452_ _4673_/B _4874_/A _3592_/D _4643_/C vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__and4_1
X_6240_ _6240_/A vssd1 vssd1 vccd1 vccd1 _6398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3383_ _4643_/C vssd1 vssd1 vccd1 vccd1 _3430_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6489__71 vssd1 vssd1 vccd1 vccd1 _6489__71/HI _6597_/A sky130_fd_sc_hd__conb_1
X_6171_ _6371_/Q _6183_/B vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__and2_1
X_5122_ _5122_/A _5168_/B vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__nand2_2
XFILLER_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5088_/A _5053_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__nor2_1
X_4004_ _4004_/A _4004_/B vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__xor2_4
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5955_ _5851_/X _5909_/X _5954_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _6322_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _5313_/A _5369_/A _5368_/A vssd1 vssd1 vccd1 vccd1 _5275_/B sky130_fd_sc_hd__and3_1
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5886_ _6421_/Q _5873_/X _5885_/X _6422_/Q vssd1 vssd1 vccd1 vccd1 _5886_/X sky130_fd_sc_hd__o22a_1
X_4837_ _4837_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4838_/C sky130_fd_sc_hd__xnor2_1
X_4768_ _4768_/A _4768_/B _4768_/C vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__and3_1
X_4699_ _4699_/A _4699_/B vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__nor2_1
X_3719_ _3720_/A _3720_/B _3741_/A vssd1 vssd1 vccd1 vccd1 _3729_/A sky130_fd_sc_hd__a21o_1
X_6369_ _6388_/CLK _6369_/D vssd1 vssd1 vccd1 vccd1 _6369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5740_ _5796_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5803_/B sky130_fd_sc_hd__or2b_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5671_/A _5665_/X vssd1 vssd1 vccd1 vccd1 _5672_/B sky130_fd_sc_hd__or2b_1
X_4622_ _5871_/B _5817_/A _5871_/A vssd1 vssd1 vccd1 vccd1 _5868_/B sky130_fd_sc_hd__o21a_2
X_4553_ _4553_/A _4553_/B vssd1 vssd1 vccd1 vccd1 _4555_/B sky130_fd_sc_hd__nor2_1
X_3504_ _3502_/A _3544_/A _3551_/A vssd1 vssd1 vccd1 vccd1 _3511_/B sky130_fd_sc_hd__a21bo_1
X_4484_ _4498_/A _4484_/B vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__xnor2_4
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3435_ _3395_/A _3466_/B _3466_/C vssd1 vssd1 vccd1 vccd1 _3467_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6223_ _6384_/Q _6387_/Q _6223_/C vssd1 vssd1 vccd1 vccd1 _6223_/X sky130_fd_sc_hd__and3_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3366_ _4307_/A vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__clkbuf_2
X_6154_ _6362_/Q _6361_/Q _6364_/Q _6363_/Q vssd1 vssd1 vccd1 vccd1 _6155_/C sky130_fd_sc_hd__or4_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5105_/A _5105_/B vssd1 vssd1 vccd1 vccd1 _5112_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3297_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3297_/Y sky130_fd_sc_hd__inv_2
X_6085_ _6099_/A _6085_/B vssd1 vssd1 vccd1 vccd1 _6085_/Y sky130_fd_sc_hd__nand2_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5048_/A _5036_/B vssd1 vssd1 vccd1 vccd1 _5038_/B sky130_fd_sc_hd__nor2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5938_ _5938_/A _5938_/B vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__nand2_1
X_5869_ _5807_/A _5867_/X _5870_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6459__41 vssd1 vssd1 vccd1 vccd1 _6459__41/HI _6564_/A sky130_fd_sc_hd__conb_1
X_3220_ _3222_/A vssd1 vssd1 vccd1 vccd1 _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3984_ _5514_/A vssd1 vssd1 vccd1 vccd1 _5425_/A sky130_fd_sc_hd__buf_2
X_5723_ _5723_/A _5723_/B vssd1 vssd1 vccd1 vccd1 _5723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5654_ _5654_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5758_/A sky130_fd_sc_hd__xor2_4
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4605_ _4593_/X _4599_/X _4602_/X _4603_/Y _4604_/X vssd1 vssd1 vccd1 vccd1 _4607_/B
+ sky130_fd_sc_hd__a32o_1
X_5585_ _5265_/Y _5269_/Y _5225_/B _5229_/X vssd1 vssd1 vccd1 vccd1 _5585_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4536_ _5672_/A _4601_/A _4536_/C vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__nand3_1
X_4467_ _4159_/Y _4167_/A _4127_/B _4129_/X vssd1 vssd1 vccd1 vccd1 _4467_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3418_ _4924_/A vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__clkbuf_4
X_4398_ _4390_/A _4396_/Y _4397_/Y vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__o21a_2
X_6206_ _6206_/A vssd1 vssd1 vccd1 vccd1 _6384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3349_ _5296_/A vssd1 vssd1 vccd1 vccd1 _5211_/A sky130_fd_sc_hd__clkbuf_2
X_6137_ _6357_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6138_/A sky130_fd_sc_hd__and2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6068_ _6060_/A _6103_/B _6063_/Y vssd1 vssd1 vccd1 vccd1 _6068_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5019_ _5019_/A _5029_/C vssd1 vssd1 vccd1 vccd1 _5020_/B sky130_fd_sc_hd__xor2_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _5487_/B vssd1 vssd1 vccd1 vccd1 _5533_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _4321_/A _4321_/B vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__nor2_2
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4252_ _5456_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4297_/A sky130_fd_sc_hd__nand3_2
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4183_ _5371_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4183_/X sky130_fd_sc_hd__and2_1
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _3960_/Y _4016_/A _3966_/Y vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5706_ _5706_/A _5706_/B vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__or2_1
X_3898_ _3898_/A _3943_/A vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__nor2_1
X_5637_ _5796_/A _5688_/A vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__or2_1
X_5568_ _5568_/A _5568_/B vssd1 vssd1 vccd1 vccd1 _5568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4519_ _4519_/A _4519_/B vssd1 vssd1 vccd1 vccd1 _4562_/A sky130_fd_sc_hd__xnor2_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5499_ _5407_/A _5545_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5500_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6429__11 vssd1 vssd1 vccd1 vccd1 _6429__11/HI _6534_/A sky130_fd_sc_hd__conb_1
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4870_ _4851_/B _4862_/A _4851_/A vssd1 vssd1 vccd1 vccd1 _4871_/B sky130_fd_sc_hd__a21oi_1
X_3821_ _5017_/A _4079_/B vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__nand2_1
X_6540_ _6540_/A _3221_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _4905_/A _4957_/B _3589_/A _4956_/A vssd1 vssd1 vccd1 vccd1 _4184_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3683_ _3683_/A _3683_/B _3703_/B vssd1 vssd1 vccd1 vccd1 _3705_/B sky130_fd_sc_hd__nand3_1
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__xnor2_2
X_5353_ _5353_/A _5353_/B _5353_/C vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__nand3_2
X_4304_ _4304_/A _4304_/B vssd1 vssd1 vccd1 vccd1 _4305_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5284_ _5311_/A _5311_/B vssd1 vssd1 vccd1 vccd1 _5326_/A sky130_fd_sc_hd__or2_1
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4235_ _4307_/A _4406_/B _4235_/C vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__and3_1
X_4166_ _4159_/Y _4162_/X _4160_/Y _4161_/Y vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__a211o_1
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _5287_/A _4221_/B vssd1 vssd1 vccd1 vccd1 _4098_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4999_ _5060_/A _5101_/B vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__and2_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6513__95 vssd1 vssd1 vccd1 vccd1 _6513__95/HI _6621_/A sky130_fd_sc_hd__conb_1
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6520__102 vssd1 vssd1 vccd1 vccd1 _6520__102/HI _6628_/A sky130_fd_sc_hd__conb_1
XFILLER_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _5248_/A _4152_/B _4021_/C vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__a21oi_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5971_ _6374_/Q _6383_/Q vssd1 vssd1 vccd1 vccd1 _5971_/X sky130_fd_sc_hd__and2b_1
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4922_ _4948_/A _4967_/B _4948_/C _4971_/B _4921_/X vssd1 vssd1 vccd1 vccd1 _4974_/B
+ sky130_fd_sc_hd__a41oi_4
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4853_ _4852_/A _4852_/B _4871_/A vssd1 vssd1 vccd1 vccd1 _4858_/B sky130_fd_sc_hd__o21bai_1
X_3804_ _3771_/Y _3804_/B vssd1 vssd1 vccd1 vccd1 _3805_/A sky130_fd_sc_hd__and2b_1
X_4784_ _4812_/B vssd1 vssd1 vccd1 vccd1 _4924_/B sky130_fd_sc_hd__clkbuf_2
X_3735_ _3735_/A _3735_/B _3735_/C vssd1 vssd1 vccd1 vccd1 _3736_/B sky130_fd_sc_hd__and3_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _5471_/B vssd1 vssd1 vccd1 vccd1 _5545_/B sky130_fd_sc_hd__clkbuf_2
X_3666_ _3669_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__nand2_1
X_3597_ _3596_/A _3597_/B vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__and2b_1
X_6385_ _6388_/CLK _6385_/D vssd1 vssd1 vccd1 vccd1 _6385_/Q sky130_fd_sc_hd__dfxtp_1
X_5336_ _5335_/A _5335_/B _5335_/C vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5267_ _5267_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__nand2_1
X_4218_ _4218_/A _4218_/B vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5198_ _5198_/A _5248_/D vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4149_ _4149_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__xor2_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _3520_/A _3520_/B vssd1 vssd1 vccd1 vccd1 _3558_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3451_ _4830_/B vssd1 vssd1 vccd1 vccd1 _4874_/A sky130_fd_sc_hd__clkbuf_2
X_6170_ _6170_/A vssd1 vssd1 vccd1 vccd1 _6371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3382_ _3538_/C vssd1 vssd1 vccd1 vccd1 _4643_/C sky130_fd_sc_hd__buf_2
X_5121_ _5121_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5052_ _5088_/A _5053_/B vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__and2_1
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4003_ _4003_/A _4003_/B vssd1 vssd1 vccd1 vccd1 _4004_/B sky130_fd_sc_hd__nor2_2
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5954_ _5954_/A _5954_/B vssd1 vssd1 vccd1 vccd1 _5954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4905_ _4905_/A _4956_/B _4905_/C vssd1 vssd1 vccd1 vccd1 _5368_/A sky130_fd_sc_hd__and3_1
X_5885_ _5936_/A _5870_/X _5884_/X _4634_/X vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4836_ _4842_/A _4842_/B vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__xor2_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4767_ _4776_/A _4754_/B _4754_/C vssd1 vssd1 vccd1 vccd1 _4768_/C sky130_fd_sc_hd__o21ai_1
X_4698_ _4697_/A _4891_/C _4749_/B _4711_/B vssd1 vssd1 vccd1 vccd1 _4699_/B sky130_fd_sc_hd__a22oi_1
X_3718_ _4855_/A _4895_/B _3718_/C _3718_/D vssd1 vssd1 vccd1 vccd1 _3741_/A sky130_fd_sc_hd__and4_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3649_ _3649_/A _3682_/A vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__nand2_1
X_6368_ _6388_/CLK _6368_/D vssd1 vssd1 vccd1 vccd1 _6368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5319_ _5364_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5365_/A sky130_fd_sc_hd__or2_1
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6299_ _6299_/A _6299_/B _6303_/C vssd1 vssd1 vccd1 vccd1 _6420_/D sky130_fd_sc_hd__nor3_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5726_/B _5668_/X _5726_/A vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4621_ _5815_/A vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4552_ _4552_/A _4552_/B _4560_/A vssd1 vssd1 vccd1 vccd1 _4553_/B sky130_fd_sc_hd__and3_1
X_3503_ _3550_/A _3550_/B vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__nand2_1
X_4483_ _3888_/X _4486_/B _4485_/A vssd1 vssd1 vccd1 vccd1 _4484_/B sky130_fd_sc_hd__a21oi_2
X_3434_ _3434_/A _3449_/A vssd1 vssd1 vccd1 vccd1 _3466_/C sky130_fd_sc_hd__xnor2_1
X_6222_ _6389_/Q _6388_/Q _6391_/Q _6390_/Q vssd1 vssd1 vccd1 vccd1 _6223_/C sky130_fd_sc_hd__and4_1
X_3365_ _6321_/Q vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6153_ _6358_/Q _6357_/Q _6360_/Q _6359_/Q vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__and4_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3296_/Y sky130_fd_sc_hd__inv_2
X_5104_ _5061_/A _5110_/A _5103_/Y vssd1 vssd1 vccd1 vccd1 _5105_/B sky130_fd_sc_hd__o21bai_1
X_6084_ _6083_/A _6083_/B _6083_/C vssd1 vssd1 vccd1 vccd1 _6085_/B sky130_fd_sc_hd__a21o_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5035_/A _5035_/B _5035_/C vssd1 vssd1 vccd1 vccd1 _5036_/B sky130_fd_sc_hd__nor3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5937_ _5937_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5938_/B sky130_fd_sc_hd__or2_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868_ _5868_/A _5868_/B _5868_/C vssd1 vssd1 vccd1 vccd1 _5870_/A sky130_fd_sc_hd__or3_2
X_4819_ _4822_/B _4822_/A vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__or2b_1
X_5799_ _4639_/A _5796_/Y _5798_/X _5751_/Y vssd1 vssd1 vccd1 vccd1 _5799_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6474__56 vssd1 vssd1 vccd1 vccd1 _6474__56/HI _6582_/A sky130_fd_sc_hd__conb_1
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5722_ _5691_/Y _5696_/X _5721_/X vssd1 vssd1 vccd1 vccd1 _5722_/X sky130_fd_sc_hd__o21a_1
X_3983_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5653_ _5766_/A _5709_/A vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__nand2_1
X_5584_ _5630_/A _5630_/B _5626_/B _5583_/Y vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__a211o_2
X_4604_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4604_/X sky130_fd_sc_hd__and2_1
X_4535_ _4535_/A _4535_/B _4535_/C vssd1 vssd1 vccd1 vccd1 _4536_/C sky130_fd_sc_hd__nand3_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4466_ _4521_/A _4521_/B _4465_/X vssd1 vssd1 vccd1 vccd1 _4515_/B sky130_fd_sc_hd__a21o_2
XFILLER_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3417_ _4780_/A vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4397_ _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4397_/Y sky130_fd_sc_hd__nand2_1
X_6205_ _6228_/A input7/X vssd1 vssd1 vccd1 vccd1 _6206_/A sky130_fd_sc_hd__and2_1
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3348_ _5356_/A vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__buf_2
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6136_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6145_/B sky130_fd_sc_hd__clkbuf_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3279_ _3279_/A vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__clkbuf_16
X_6067_ _6074_/B vssd1 vssd1 vccd1 vccd1 _6103_/B sky130_fd_sc_hd__clkbuf_2
X_5018_ _5018_/A _5031_/A vssd1 vssd1 vccd1 vccd1 _5029_/C sky130_fd_sc_hd__xnor2_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4320_ _4349_/A _4349_/B vssd1 vssd1 vccd1 vccd1 _4321_/B sky130_fd_sc_hd__and2b_1
X_4251_ _4251_/A _4251_/B vssd1 vssd1 vccd1 vccd1 _4463_/B sky130_fd_sc_hd__xnor2_2
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4182_ _4182_/A _4182_/B vssd1 vssd1 vccd1 vccd1 _4194_/A sky130_fd_sc_hd__or2_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3966_ _3966_/A _3966_/B vssd1 vssd1 vccd1 vccd1 _3966_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5705_ _5712_/A _5560_/B _5560_/C vssd1 vssd1 vccd1 vccd1 _5706_/B sky130_fd_sc_hd__a21oi_1
X_3897_ _3960_/A _4008_/B vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__nand2_1
X_5636_ _5636_/A _5636_/B vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__xnor2_4
X_5567_ _5565_/A _5565_/B _5680_/A vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__o21bai_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5498_ _5498_/A _5498_/B vssd1 vssd1 vccd1 vccd1 _5517_/A sky130_fd_sc_hd__xor2_2
X_4518_ _5805_/A _4547_/A vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__xnor2_1
X_4449_ _4544_/B _4449_/B vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__or2_1
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6119_ _6119_/A vssd1 vssd1 vccd1 vccd1 _6351_/D sky130_fd_sc_hd__clkbuf_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6444__26 vssd1 vssd1 vccd1 vccd1 _6444__26/HI _6549_/A sky130_fd_sc_hd__conb_1
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _3903_/B vssd1 vssd1 vccd1 vccd1 _4079_/B sky130_fd_sc_hd__buf_2
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3751_ _4872_/A vssd1 vssd1 vccd1 vccd1 _4956_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3682_ _3682_/A _3682_/B _3682_/C vssd1 vssd1 vccd1 vccd1 _3690_/C sky130_fd_sc_hd__and3_1
X_5421_ _5421_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5640_/A sky130_fd_sc_hd__xnor2_4
X_5352_ _5324_/A _5196_/B _5349_/X _5351_/Y vssd1 vssd1 vccd1 vccd1 _5353_/C sky130_fd_sc_hd__a31o_1
XFILLER_114_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4303_ _5246_/A _4347_/B _4301_/A _4302_/X vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__a31o_2
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5283_ _5283_/A _5283_/B vssd1 vssd1 vccd1 vccd1 _5311_/B sky130_fd_sc_hd__xor2_1
X_4234_ _4236_/A _4234_/B vssd1 vssd1 vccd1 vccd1 _4235_/C sky130_fd_sc_hd__nor2_1
XFILLER_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4165_ _4509_/A vssd1 vssd1 vccd1 vccd1 _4165_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4096_/A _4096_/B vssd1 vssd1 vccd1 vccd1 _4114_/C sky130_fd_sc_hd__nor2_1
XFILLER_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4998_ _5335_/B vssd1 vssd1 vccd1 vccd1 _5101_/B sky130_fd_sc_hd__buf_2
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3949_ _3947_/A _3947_/B _3981_/A vssd1 vssd1 vccd1 vccd1 _3949_/X sky130_fd_sc_hd__a21bo_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6599_ _6599_/A _3294_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
X_5619_ _5619_/A _5619_/B _5619_/C vssd1 vssd1 vccd1 vccd1 _5666_/B sky130_fd_sc_hd__nand3_2
XFILLER_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _6383_/Q _6374_/Q vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__and2b_1
X_4921_ _4970_/A _4793_/X _4970_/B vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__o21a_1
X_4852_ _4852_/A _4852_/B _4871_/A vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__or3b_1
X_3803_ _3818_/A vssd1 vssd1 vccd1 vccd1 _5684_/A sky130_fd_sc_hd__buf_2
X_4783_ _4787_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _4794_/B sky130_fd_sc_hd__and2_1
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3734_ _3732_/A _3731_/C _3731_/B vssd1 vssd1 vccd1 vccd1 _3757_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3665_ _3669_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__or2_1
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5404_ _5510_/B vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__clkbuf_2
X_3596_ _3596_/A _3597_/B vssd1 vssd1 vccd1 vccd1 _3637_/B sky130_fd_sc_hd__xor2_1
X_6384_ _6388_/CLK _6384_/D vssd1 vssd1 vccd1 vccd1 _6384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5335_ _5335_/A _5335_/B _5335_/C vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__and3_1
X_5266_ _5266_/A _5258_/A vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__or2b_1
X_4217_ _5324_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4218_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5197_ _5000_/A _5240_/B _5233_/A _5242_/A vssd1 vssd1 vccd1 vccd1 _5201_/B sky130_fd_sc_hd__a31oi_1
XFILLER_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4111_/X _4148_/B vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__and2b_1
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4079_ _5214_/A _4079_/B _4079_/C _4079_/D vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__and4_2
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3450_ _6328_/Q vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__buf_2
X_3381_ _3409_/A _3409_/B _6343_/Q vssd1 vssd1 vccd1 vccd1 _3538_/C sky130_fd_sc_hd__a21o_1
X_5120_ _5120_/A _5132_/B vssd1 vssd1 vccd1 vccd1 _5126_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5606_/A _5606_/B vssd1 vssd1 vccd1 vccd1 _5053_/B sky130_fd_sc_hd__xnor2_1
X_4002_ _4005_/A _4005_/B _4005_/C vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__and3_1
X_6527__109 vssd1 vssd1 vccd1 vccd1 _6527__109/HI _6635_/A sky130_fd_sc_hd__conb_1
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _5953_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__xnor2_1
X_4904_ _4904_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__xor2_2
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5884_ _5866_/X _5796_/Y _5798_/X _5871_/X vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4835_ _4891_/A _4854_/B vssd1 vssd1 vccd1 vccd1 _4842_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _4770_/B _4760_/X _4810_/B _4765_/X vssd1 vssd1 vccd1 vccd1 _4768_/B sky130_fd_sc_hd__a31o_1
X_3717_ _4850_/A _3718_/C _3716_/D _4830_/A vssd1 vssd1 vccd1 vccd1 _3720_/B sky130_fd_sc_hd__a22o_1
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4697_ _4697_/A _4697_/B _4891_/C _4749_/B vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__and4_1
X_3648_ _3649_/A _3648_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3682_/A sky130_fd_sc_hd__nand3_2
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6367_ _6388_/CLK _6367_/D vssd1 vssd1 vccd1 vccd1 _6367_/Q sky130_fd_sc_hd__dfxtp_1
X_3579_ _3409_/A _3359_/A _6040_/A vssd1 vssd1 vccd1 vccd1 _3671_/B sky130_fd_sc_hd__a21o_2
XFILLER_115_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5318_ _5318_/A _5318_/B vssd1 vssd1 vccd1 vccd1 _5364_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6298_ _6420_/Q _6298_/B _6418_/Q vssd1 vssd1 vccd1 vccd1 _6303_/C sky130_fd_sc_hd__and3_1
X_5249_ _5249_/A _5249_/B vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _6344_/Q vssd1 vssd1 vccd1 vccd1 _5817_/A sky130_fd_sc_hd__clkbuf_2
X_4551_ _5015_/A vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__clkbuf_4
X_3502_ _3502_/A _3502_/B vssd1 vssd1 vccd1 vccd1 _3550_/B sky130_fd_sc_hd__xnor2_1
X_4482_ _4482_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__and2_1
X_3433_ _3592_/C vssd1 vssd1 vccd1 vccd1 _3466_/B sky130_fd_sc_hd__clkbuf_2
X_6221_ _6221_/A vssd1 vssd1 vccd1 vccd1 _6391_/D sky130_fd_sc_hd__clkbuf_1
X_6152_ _6362_/Q _6361_/Q _6364_/Q _6363_/Q vssd1 vssd1 vccd1 vccd1 _6152_/X sky130_fd_sc_hd__and4_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5103_ _4989_/A _5353_/B _5128_/B _3960_/A vssd1 vssd1 vccd1 vccd1 _5103_/Y sky130_fd_sc_hd__a22oi_2
X_3364_ _3364_/A _3364_/B vssd1 vssd1 vccd1 vccd1 _5745_/B sky130_fd_sc_hd__nand2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3295_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6083_ _6083_/A _6083_/B _6083_/C vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__and3_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5034_ _5035_/A _5035_/B _5035_/C vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__o21a_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5936_ _5936_/A _5944_/A vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5867_ _5758_/Y _5866_/X _5823_/C _5759_/Y vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__a22o_1
X_4818_ _4811_/A _4811_/B _4817_/X vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__a21o_1
X_5798_ _5805_/B _5797_/X vssd1 vssd1 vccd1 vccd1 _5798_/X sky130_fd_sc_hd__or2b_1
X_4749_ _4888_/A _4749_/B vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6419_ _6423_/CLK _6419_/D vssd1 vssd1 vccd1 vccd1 _6419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3982_ _6317_/Q vssd1 vssd1 vccd1 vccd1 _5518_/A sky130_fd_sc_hd__clkbuf_2
X_5721_ _5691_/Y _5696_/X _5716_/Y _5719_/Y _5720_/Y vssd1 vssd1 vccd1 vccd1 _5721_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5652_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5709_/A sky130_fd_sc_hd__xor2_4
X_5583_ _5583_/A _5583_/B vssd1 vssd1 vccd1 vccd1 _5583_/Y sky130_fd_sc_hd__nor2_1
X_4603_ _4602_/A _4602_/B _4598_/X vssd1 vssd1 vccd1 vccd1 _4603_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4534_ _4535_/A _4535_/B _4535_/C vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__a21o_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4465_ _4250_/B _4465_/B vssd1 vssd1 vccd1 vccd1 _4465_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4396_ _5324_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4396_/Y sky130_fd_sc_hd__nand2_1
X_3416_ _4651_/A vssd1 vssd1 vccd1 vccd1 _4780_/A sky130_fd_sc_hd__buf_2
X_6204_ _5911_/X _6199_/X _6200_/X _6203_/X _6335_/D vssd1 vssd1 vccd1 vccd1 _6383_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3347_ _5433_/A vssd1 vssd1 vccd1 vccd1 _5356_/A sky130_fd_sc_hd__buf_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _6135_/A vssd1 vssd1 vccd1 vccd1 _6357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6066_ _6341_/Q _6074_/B vssd1 vssd1 vccd1 vccd1 _6077_/B sky130_fd_sc_hd__xor2_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5017_ _5017_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5031_/A sky130_fd_sc_hd__and2_1
X_3278_ _3278_/A vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5919_ _5954_/A _5919_/B vssd1 vssd1 vccd1 vccd1 _5919_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4465_/B _4250_/B vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__xnor2_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4181_ _4109_/A _4212_/B _4136_/C vssd1 vssd1 vccd1 vccd1 _4182_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3965_ _5282_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__nand2_1
X_3896_ _4263_/B vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5704_ _5761_/A _5704_/B vssd1 vssd1 vccd1 vccd1 _5704_/Y sky130_fd_sc_hd__xnor2_1
X_5635_ _5629_/Y _5633_/Y _5634_/X vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__a21o_1
X_5566_ _5679_/B _5686_/A _5565_/X vssd1 vssd1 vccd1 vccd1 _5680_/A sky130_fd_sc_hd__a21boi_1
X_5497_ _5497_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__xor2_2
X_4517_ _5750_/A _4540_/A vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__xor2_1
X_4448_ _4448_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4449_/B sky130_fd_sc_hd__and2_1
X_4379_ _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__or2_1
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6118_ _6350_/Q _6314_/B vssd1 vssd1 vccd1 vccd1 _6119_/A sky130_fd_sc_hd__and2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6049_ _6049_/A _6049_/B vssd1 vssd1 vccd1 vccd1 _6050_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3750_ _4872_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _4957_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3681_ _3681_/A _3681_/B vssd1 vssd1 vccd1 vccd1 _3694_/B sky130_fd_sc_hd__xor2_2
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5420_ _5422_/A _5422_/B _5419_/X vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5351_ _5351_/A _5351_/B vssd1 vssd1 vccd1 vccd1 _5351_/Y sky130_fd_sc_hd__nor2_1
X_4302_ _5353_/A _4302_/B _4318_/A vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__and3_1
X_5282_ _5282_/A _5458_/B vssd1 vssd1 vccd1 vccd1 _5283_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _5441_/A _4387_/B _4336_/A _4272_/A vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__a22oi_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4164_ _4127_/B _4129_/X _4159_/Y _4167_/A vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__o211ai_2
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4095_ _4095_/A _4263_/B _4095_/C vssd1 vssd1 vccd1 vccd1 _4096_/B sky130_fd_sc_hd__and3_1
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4997_ _5257_/B vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3948_ _3948_/A _3948_/B _3948_/C vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__nand3_1
X_3879_ _3878_/B _3879_/B vssd1 vssd1 vccd1 vccd1 _3879_/X sky130_fd_sc_hd__and2b_1
X_6598_ _6598_/A _3293_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
X_5618_ _5619_/A _5619_/B _5619_/C vssd1 vssd1 vccd1 vccd1 _5666_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5549_ _5549_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__nor2_2
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6423_/CLK
+ sky130_fd_sc_hd__clkbuf_2
X_6504__86 vssd1 vssd1 vccd1 vccd1 _6504__86/HI _6612_/A sky130_fd_sc_hd__conb_1
XFILLER_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _4970_/A _4970_/B vssd1 vssd1 vccd1 vccd1 _4971_/B sky130_fd_sc_hd__or2_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4851_ _4851_/A _4851_/B _4862_/A vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__and3_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ _3843_/B _3802_/B vssd1 vssd1 vccd1 vccd1 _3812_/A sky130_fd_sc_hd__or2_1
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__xor2_1
X_3733_ _3759_/A _3759_/B _3759_/C vssd1 vssd1 vccd1 vccd1 _3733_/X sky130_fd_sc_hd__a21o_1
X_3664_ _3681_/A _3681_/B _3663_/X vssd1 vssd1 vccd1 vccd1 _3669_/B sky130_fd_sc_hd__o21ai_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5403_ _5368_/B _5403_/B vssd1 vssd1 vccd1 vccd1 _5510_/B sky130_fd_sc_hd__and2b_1
X_3595_ _3626_/A _3626_/B _3594_/X vssd1 vssd1 vccd1 vccd1 _3597_/B sky130_fd_sc_hd__a21bo_1
X_6383_ _6388_/CLK _6383_/D vssd1 vssd1 vccd1 vccd1 _6383_/Q sky130_fd_sc_hd__dfxtp_1
X_5334_ _5290_/A _5248_/D _5325_/A _5333_/Y vssd1 vssd1 vccd1 vccd1 _5335_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5265_ _5268_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5265_/Y sky130_fd_sc_hd__nand2_1
X_4216_ _4237_/A _4237_/B _4213_/X vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__o21ba_1
X_5196_ _5198_/A _5196_/B _5196_/C vssd1 vssd1 vccd1 vccd1 _5242_/A sky130_fd_sc_hd__and3_1
XFILLER_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4147_ _4144_/A _4144_/B _4145_/B _4146_/Y vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__o31a_1
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _5168_/A _3818_/B _4069_/B _4076_/X vssd1 vssd1 vccd1 vccd1 _4079_/D sky130_fd_sc_hd__a211o_1
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3380_ _3466_/A vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5050_ _5601_/A _5050_/B vssd1 vssd1 vccd1 vccd1 _5606_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4001_ _3997_/X _3998_/Y _3980_/Y _3996_/X vssd1 vssd1 vccd1 vccd1 _4005_/C sky130_fd_sc_hd__o211ai_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5952_ _5945_/A _5950_/B _5951_/X vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4903_ _4955_/B _4903_/B vssd1 vssd1 vccd1 vccd1 _5313_/A sky130_fd_sc_hd__nor2_1
XFILLER_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5883_ _6420_/Q _5869_/Y _5873_/X _6421_/Q _5882_/X vssd1 vssd1 vccd1 vccd1 _5883_/X
+ sky130_fd_sc_hd__a221o_1
X_4834_ _4872_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4837_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4765_ _4764_/A _4891_/D _4828_/A _4765_/D vssd1 vssd1 vccd1 vccd1 _4765_/X sky130_fd_sc_hd__and4b_1
X_3716_ _4800_/A _4874_/A _3716_/C _3716_/D vssd1 vssd1 vccd1 vccd1 _3720_/A sky130_fd_sc_hd__nand4_1
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4696_ _4728_/A _4854_/B vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3647_/A _3718_/C vssd1 vssd1 vccd1 vccd1 _3648_/C sky130_fd_sc_hd__nand2_1
X_6366_ _6388_/CLK _6366_/D vssd1 vssd1 vccd1 vccd1 _6366_/Q sky130_fd_sc_hd__dfxtp_1
X_3578_ _6336_/Q vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5317_ _5317_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5364_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6297_ _6298_/B _6294_/A _6420_/Q vssd1 vssd1 vccd1 vccd1 _6299_/B sky130_fd_sc_hd__a21oi_1
X_5248_ _5248_/A _5248_/B _5290_/B _5248_/D vssd1 vssd1 vccd1 vccd1 _5249_/B sky130_fd_sc_hd__and4_1
X_6495__77 vssd1 vssd1 vccd1 vccd1 _6495__77/HI _6603_/A sky130_fd_sc_hd__conb_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5179_ _5178_/A _5212_/A _5170_/X _5121_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5182_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _5684_/A _4550_/B vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__xor2_1
X_3501_ _3506_/A _3501_/B vssd1 vssd1 vccd1 vccd1 _3550_/A sky130_fd_sc_hd__xnor2_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4481_ _4488_/A _4488_/B _4488_/C _3928_/A vssd1 vssd1 vccd1 vccd1 _4486_/B sky130_fd_sc_hd__a31o_2
X_6220_ _6390_/Q _6232_/B vssd1 vssd1 vccd1 vccd1 _6221_/A sky130_fd_sc_hd__and2_1
X_3432_ _3628_/C vssd1 vssd1 vccd1 vccd1 _3592_/C sky130_fd_sc_hd__clkbuf_4
X_6151_ _6151_/A vssd1 vssd1 vccd1 vccd1 _6364_/D sky130_fd_sc_hd__clkbuf_1
X_3363_ _5871_/B _6344_/Q _5815_/A vssd1 vssd1 vccd1 vccd1 _3364_/B sky130_fd_sc_hd__or3b_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5102_ _5102_/A _5248_/D vssd1 vssd1 vccd1 vccd1 _5110_/A sky130_fd_sc_hd__nand2_2
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3294_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3294_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6082_ _6343_/Q _6088_/B vssd1 vssd1 vccd1 vccd1 _6083_/C sky130_fd_sc_hd__xor2_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5033_ _5045_/B _5033_/B vssd1 vssd1 vccd1 vccd1 _5035_/C sky130_fd_sc_hd__and2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5935_ _5785_/X _5933_/X _5934_/Y vssd1 vssd1 vccd1 vccd1 _6319_/D sky130_fd_sc_hd__o21a_1
X_5866_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4817_ _4826_/A _4826_/B vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__and2b_1
X_5797_ _5789_/A _4617_/C _5789_/B _4617_/B vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__a31o_1
X_4748_ _4747_/A _4747_/B _4747_/C vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__a21oi_1
X_4679_ _4679_/A _4679_/B vssd1 vssd1 vccd1 vccd1 _4680_/B sky130_fd_sc_hd__xnor2_1
X_6418_ _6423_/CLK _6418_/D vssd1 vssd1 vccd1 vccd1 _6418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6349_ _6401_/CLK _6349_/D vssd1 vssd1 vccd1 vccd1 _6349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3981_ _3981_/A _3981_/B _3981_/C vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__and3_1
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5720_ _5720_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _5669_/A vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__clkbuf_2
X_5582_ _5625_/B _5625_/C _5625_/A vssd1 vssd1 vccd1 vccd1 _5626_/B sky130_fd_sc_hd__a21oi_1
X_4602_ _4602_/A _4602_/B vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__xor2_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4533_ _4533_/A _4533_/B vssd1 vssd1 vccd1 vccd1 _4535_/C sky130_fd_sc_hd__xnor2_4
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4464_ _4519_/A _4519_/B _4463_/X vssd1 vssd1 vccd1 vccd1 _4521_/B sky130_fd_sc_hd__a21o_2
X_6203_ _6377_/Q _6203_/B _6203_/C vssd1 vssd1 vccd1 vccd1 _6203_/X sky130_fd_sc_hd__or3_1
X_4395_ _4411_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__or2_2
X_3415_ _4756_/A vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3346_ _4014_/A vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__clkbuf_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6134_/A input4/X vssd1 vssd1 vccd1 vccd1 _6135_/A sky130_fd_sc_hd__and2_1
X_6465__47 vssd1 vssd1 vccd1 vccd1 _6465__47/HI _6570_/A sky130_fd_sc_hd__conb_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6060_/A _6036_/X _6064_/X _6015_/X vssd1 vssd1 vccd1 vccd1 _6340_/D sky130_fd_sc_hd__o211a_1
X_5016_ _5030_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__nand2_1
X_3277_ _3278_/A vssd1 vssd1 vccd1 vccd1 _3277_/Y sky130_fd_sc_hd__inv_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5918_ _5918_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5919_/B sky130_fd_sc_hd__xnor2_1
X_5849_ _6106_/A _6104_/A _6104_/B vssd1 vssd1 vccd1 vccd1 _5849_/X sky130_fd_sc_hd__or3_1
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4180_ _4180_/A _4180_/B vssd1 vssd1 vccd1 vccd1 _4223_/A sky130_fd_sc_hd__xor2_1
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3964_ _4169_/C vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3895_ _4066_/B vssd1 vssd1 vccd1 vccd1 _4263_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5703_ _5703_/A _5703_/B vssd1 vssd1 vccd1 vccd1 _5704_/B sky130_fd_sc_hd__nor2_1
X_5634_ _5634_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5634_/X sky130_fd_sc_hd__xor2_1
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5565_ _5565_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _5565_/X sky130_fd_sc_hd__xor2_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5496_ _5509_/A _5496_/B vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__or2_1
X_4516_ _5805_/A _4547_/A vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__nand2_1
X_4447_ _4567_/A _4559_/B vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__or2_1
X_4378_ _4380_/A _4380_/B _4377_/X vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__a21o_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6314_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3329_ _3333_/A vssd1 vssd1 vccd1 vccd1 _3329_/Y sky130_fd_sc_hd__inv_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _6038_/A _6059_/A _6039_/X vssd1 vssd1 vccd1 vccd1 _6049_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3680_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5350_ _5350_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _5351_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4301_ _4301_/A _4301_/B vssd1 vssd1 vccd1 vccd1 _4318_/A sky130_fd_sc_hd__xnor2_2
X_5281_ _5281_/A _5350_/B vssd1 vssd1 vccd1 vccd1 _5311_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4232_ _4383_/C vssd1 vssd1 vccd1 vccd1 _4336_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ _4160_/Y _4161_/Y _4159_/Y _4162_/X vssd1 vssd1 vccd1 vccd1 _4167_/A sky130_fd_sc_hd__o211ai_4
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4094_ _5288_/A _4008_/B _4095_/C vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__a21oi_1
X_6435__17 vssd1 vssd1 vccd1 vccd1 _6435__17/HI _6540_/A sky130_fd_sc_hd__conb_1
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4996_ _5168_/B vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__clkbuf_2
X_3947_ _3947_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _3948_/C sky130_fd_sc_hd__xor2_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3878_ _3879_/B _3878_/B vssd1 vssd1 vccd1 vccd1 _3891_/B sky130_fd_sc_hd__xnor2_1
X_5617_ _5585_/Y _5617_/B vssd1 vssd1 vccd1 vccd1 _5619_/C sky130_fd_sc_hd__and2b_1
X_6597_ _6597_/A _3291_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_5548_ _5514_/A _5555_/D _5533_/C vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__a21oi_1
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5479_ _5478_/A _5479_/B vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__and2b_1
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4850_/A _4850_/B _4874_/C vssd1 vssd1 vccd1 vccd1 _4862_/A sky130_fd_sc_hd__nand3_1
X_3801_ _3818_/A _3849_/B _3800_/C vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__a21oi_1
X_4781_ _4624_/A _4716_/X _4779_/Y _4780_/X vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__a211o_1
X_3732_ _3732_/A _3757_/A vssd1 vssd1 vccd1 vccd1 _3759_/C sky130_fd_sc_hd__nand2_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3663_ _3663_/A _3690_/A vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__or2_1
X_5402_ _4624_/A _4956_/B _4957_/A _4957_/C _4957_/B vssd1 vssd1 vccd1 vccd1 _5403_/B
+ sky130_fd_sc_hd__a221o_1
X_6382_ _6396_/CLK _6382_/D vssd1 vssd1 vccd1 vccd1 _6382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5333_ _5333_/A _5351_/A vssd1 vssd1 vccd1 vccd1 _5333_/Y sky130_fd_sc_hd__nor2_1
X_3594_ _3594_/A _3593_/B vssd1 vssd1 vccd1 vccd1 _3594_/X sky130_fd_sc_hd__or2b_1
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5264_ _5264_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _5268_/B sky130_fd_sc_hd__xnor2_2
X_4215_ _5458_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4237_/B sky130_fd_sc_hd__nand2_1
X_5195_ _5195_/A _5233_/A vssd1 vssd1 vccd1 vccd1 _5196_/C sky130_fd_sc_hd__xnor2_1
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _4178_/A _4178_/B vssd1 vssd1 vccd1 vccd1 _4146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4069_/B _4076_/X _5121_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _4079_/C sky130_fd_sc_hd__o211ai_4
XFILLER_56_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4979_ _4995_/A _4995_/B _4979_/C _4979_/D vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__or4_4
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4000_ _3980_/Y _3996_/X _3997_/X _3998_/Y vssd1 vssd1 vccd1 vccd1 _4005_/B sky130_fd_sc_hd__a211o_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _5842_/A _5944_/A _5946_/A vssd1 vssd1 vccd1 vccd1 _5951_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4902_ _4902_/A _4902_/B _4902_/C vssd1 vssd1 vccd1 vccd1 _4903_/B sky130_fd_sc_hd__nor3_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5882_ _6420_/Q _5869_/Y _5878_/X _5881_/X vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4833_ _4832_/A _4832_/B _4852_/A vssd1 vssd1 vccd1 vccd1 _4838_/B sky130_fd_sc_hd__a21o_1
X_4764_ _4764_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__xor2_2
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3715_ _3706_/A _3706_/C _3706_/B vssd1 vssd1 vccd1 vccd1 _3730_/C sky130_fd_sc_hd__a21o_1
X_4695_ _4758_/B vssd1 vssd1 vccd1 vccd1 _4854_/B sky130_fd_sc_hd__buf_2
X_3646_ _3646_/A _3672_/A _3646_/C _3699_/D vssd1 vssd1 vccd1 vccd1 _3648_/B sky130_fd_sc_hd__nand4_1
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3577_ _3577_/A _3577_/B vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__xnor2_1
X_6365_ _6396_/CLK _6365_/D vssd1 vssd1 vccd1 vccd1 _6365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5316_ _5316_/A _5514_/B vssd1 vssd1 vccd1 vccd1 _5318_/B sky130_fd_sc_hd__nand2_1
X_6296_ _6298_/B _6294_/A _6295_/Y vssd1 vssd1 vccd1 vccd1 _6419_/D sky130_fd_sc_hd__a21oi_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5247_ _3974_/A _5353_/B _5128_/B _5248_/A vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__a22oi_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5178_ _5178_/A _5212_/A vssd1 vssd1 vccd1 vccd1 _5182_/A sky130_fd_sc_hd__nor2_1
X_4129_ _4127_/A _4125_/X _4118_/C _4121_/B vssd1 vssd1 vccd1 vccd1 _4129_/X sky130_fd_sc_hd__o211a_1
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3500_ _4711_/A _3718_/D vssd1 vssd1 vccd1 vccd1 _3501_/B sky130_fd_sc_hd__nand2_1
X_4480_ _4476_/X _4479_/Y _4493_/A vssd1 vssd1 vccd1 vccd1 _4488_/C sky130_fd_sc_hd__a21o_1
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3431_ _3409_/A _3359_/A _6340_/Q vssd1 vssd1 vccd1 vccd1 _3628_/C sky130_fd_sc_hd__a21o_1
X_6150_ _6363_/Q _6164_/B vssd1 vssd1 vccd1 vccd1 _6151_/A sky130_fd_sc_hd__and2_1
X_3362_ _3409_/B vssd1 vssd1 vccd1 vccd1 _5871_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5101_ _5118_/A _5101_/B vssd1 vssd1 vccd1 vccd1 _5105_/A sky130_fd_sc_hd__nand2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3293_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3293_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6081_ _6074_/A _6032_/X _6080_/X _5948_/X vssd1 vssd1 vccd1 vccd1 _6342_/D sky130_fd_sc_hd__o211a_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5032_ _5028_/A _5214_/B _5029_/B _3818_/A vssd1 vssd1 vccd1 vccd1 _5033_/B sky130_fd_sc_hd__a22o_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5934_ _5785_/X _5933_/X _6299_/A vssd1 vssd1 vccd1 vccd1 _5934_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5865_ _5848_/A _5871_/A _6103_/A vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__and3b_1
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4816_ _4816_/A _4816_/B vssd1 vssd1 vccd1 vccd1 _4826_/B sky130_fd_sc_hd__xnor2_2
XFILLER_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5796_ _5796_/A _5796_/B vssd1 vssd1 vccd1 vccd1 _5796_/Y sky130_fd_sc_hd__xnor2_1
X_4747_ _4747_/A _4747_/B _4747_/C vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__and3_1
X_4678_ _4692_/C _4678_/B vssd1 vssd1 vccd1 vccd1 _4679_/B sky130_fd_sc_hd__xor2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6417_ _6423_/CLK _6417_/D vssd1 vssd1 vccd1 vccd1 _6417_/Q sky130_fd_sc_hd__dfxtp_1
X_3629_ _6328_/Q vssd1 vssd1 vccd1 vccd1 _3672_/A sky130_fd_sc_hd__clkbuf_2
X_6348_ _6401_/CLK _6348_/D vssd1 vssd1 vccd1 vccd1 _6348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6279_ _6413_/Q _6283_/C vssd1 vssd1 vccd1 vccd1 _6280_/B sky130_fd_sc_hd__and2_1
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _3981_/A _3981_/B _3981_/C vssd1 vssd1 vccd1 vccd1 _3980_/Y sky130_fd_sc_hd__nand3_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5650_ _5650_/A _5650_/B vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__xnor2_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4601_ _4601_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4602_/B sky130_fd_sc_hd__and2_1
X_5581_ _5636_/A _5636_/B _5580_/X vssd1 vssd1 vccd1 vccd1 _5630_/B sky130_fd_sc_hd__a21o_2
X_4532_ _5789_/A _4569_/A vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__xnor2_1
X_4463_ _4293_/B _4463_/B vssd1 vssd1 vccd1 vccd1 _4463_/X sky130_fd_sc_hd__and2b_1
X_3414_ _3421_/A _3421_/B vssd1 vssd1 vccd1 vccd1 _3441_/B sky130_fd_sc_hd__nand2_1
X_6202_ _6380_/Q _6379_/Q _6382_/Q _6381_/Q vssd1 vssd1 vccd1 vccd1 _6203_/C sky130_fd_sc_hd__or4_1
X_4394_ _4394_/A _4394_/B vssd1 vssd1 vccd1 vccd1 _4411_/B sky130_fd_sc_hd__or2_1
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3345_ _4104_/A vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__buf_2
X_6133_ _6349_/Q _6349_/D _6129_/X _6132_/X vssd1 vssd1 vccd1 vccd1 _6356_/D sky130_fd_sc_hd__a31o_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3276_ _3278_/A vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__inv_2
X_6064_ _6062_/X _6063_/Y _6036_/A vssd1 vssd1 vccd1 vccd1 _6064_/X sky130_fd_sc_hd__a21bo_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__nand2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5917_ _5915_/X _5917_/B vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__and2b_1
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5848_ _5848_/A vssd1 vssd1 vccd1 vccd1 _6104_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779_ _5779_/A _5779_/B vssd1 vssd1 vccd1 vccd1 _5779_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3963_ _4014_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__nand2_1
X_3894_ _3894_/A _3894_/B vssd1 vssd1 vccd1 vccd1 _4066_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_5702_ _5702_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _5703_/B sky130_fd_sc_hd__nor2_1
X_5633_ _5633_/A _5633_/B vssd1 vssd1 vccd1 vccd1 _5633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564_ _5693_/A _5564_/B _5699_/A vssd1 vssd1 vccd1 vccd1 _5686_/A sky130_fd_sc_hd__nand3_1
X_4515_ _4515_/A _4515_/B vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__xor2_4
X_5495_ _5493_/B _5495_/B vssd1 vssd1 vccd1 vccd1 _5496_/B sky130_fd_sc_hd__and2b_1
X_4446_ _4446_/A _4446_/B vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4377_ _4377_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__and2_1
XFILLER_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3328_ _3334_/A vssd1 vssd1 vccd1 vccd1 _3333_/A sky130_fd_sc_hd__buf_12
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A vssd1 vssd1 vccd1 vccd1 _6350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6047_ _6047_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259_ _3260_/A vssd1 vssd1 vccd1 vccd1 _3259_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4300_ _5425_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4301_/B sky130_fd_sc_hd__nand2_1
X_5280_ _5406_/A _5458_/B vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__nand2_2
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4231_ _4231_/A vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4162_ _4121_/Y _4158_/X _4150_/X _4157_/X vssd1 vssd1 vccd1 vccd1 _4162_/X sky130_fd_sc_hd__a211o_1
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4093_ _5317_/A _4140_/B vssd1 vssd1 vccd1 vccd1 _4095_/C sky130_fd_sc_hd__and2_1
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _4995_/A _4995_/B vssd1 vssd1 vccd1 vccd1 _5168_/B sky130_fd_sc_hd__xnor2_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3946_ _3933_/A _3934_/A _5068_/A _4079_/B vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3877_ _3875_/A _3898_/A _3893_/A vssd1 vssd1 vccd1 vccd1 _3878_/B sky130_fd_sc_hd__o21ba_1
X_6596_ _6596_/A _3290_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_5616_ _4274_/A _5045_/B _5614_/X _5609_/A _5615_/X vssd1 vssd1 vccd1 vccd1 _5634_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547_ _5547_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _5553_/A sky130_fd_sc_hd__xor2_2
XFILLER_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5478_ _5478_/A _5479_/B vssd1 vssd1 vccd1 vccd1 _5494_/B sky130_fd_sc_hd__xor2_1
X_4429_ _4441_/A _4408_/B _4428_/Y vssd1 vssd1 vccd1 vccd1 _4433_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4780_ _4780_/A _4891_/D _4780_/C vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__and3_1
X_3800_ _3818_/A _3849_/B _3800_/C vssd1 vssd1 vccd1 vccd1 _3843_/B sky130_fd_sc_hd__and3_1
X_3731_ _3732_/A _3731_/B _3731_/C vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__nand3_2
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3662_ _3663_/A _3690_/A vssd1 vssd1 vccd1 vccd1 _3681_/B sky130_fd_sc_hd__xnor2_2
X_3593_ _3594_/A _3593_/B vssd1 vssd1 vccd1 vccd1 _3626_/B sky130_fd_sc_hd__xnor2_2
X_5401_ _5401_/A _5401_/B vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__xor2_2
X_6381_ _6396_/CLK _6381_/D vssd1 vssd1 vccd1 vccd1 _6381_/Q sky130_fd_sc_hd__dfxtp_1
X_5332_ _5356_/A _5458_/B vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__nand2_2
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5263_ _5272_/A _5272_/B _5262_/X vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__o21ai_2
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4214_ _4211_/Y _4212_/Y _4213_/X vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__a21o_1
X_5194_ _5316_/A _5492_/B _5492_/C vssd1 vssd1 vccd1 vccd1 _5233_/A sky130_fd_sc_hd__and3_1
X_4145_ _4145_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4076_ _4069_/A _4069_/B _5095_/A _4174_/B vssd1 vssd1 vccd1 vccd1 _4076_/X sky130_fd_sc_hd__and4bb_1
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _4978_/A _4978_/B _4978_/C vssd1 vssd1 vccd1 vccd1 _4979_/D sky130_fd_sc_hd__and3_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3929_ _5154_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _3930_/C sky130_fd_sc_hd__and2_1
XFILLER_105_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6579_ _6579_/A _3269_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_117_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5950_ _5950_/A _5950_/B vssd1 vssd1 vccd1 vccd1 _5953_/A sky130_fd_sc_hd__xnor2_1
X_4901_ _4902_/B _4902_/C _4902_/A vssd1 vssd1 vccd1 vccd1 _4955_/B sky130_fd_sc_hd__o21a_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5881_ _6294_/A _5875_/X _6298_/B vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _4832_/A _4832_/B _4852_/A vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4763_ _4763_/A _4805_/C _4895_/D vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__and3_1
X_3714_ _3712_/A _3711_/C _3711_/B vssd1 vssd1 vccd1 vccd1 _3759_/B sky130_fd_sc_hd__a21o_1
X_4694_ _4694_/A _4694_/B vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__xor2_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3645_ _3672_/A _3566_/A _3570_/C _4755_/B vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__a22o_1
X_3576_ _3576_/A _3576_/B vssd1 vssd1 vccd1 vccd1 _3577_/B sky130_fd_sc_hd__or2_1
X_6364_ _6401_/CLK _6364_/D vssd1 vssd1 vccd1 vccd1 _6364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6295_ _6298_/B _6294_/A _6134_/A vssd1 vssd1 vccd1 vccd1 _6295_/Y sky130_fd_sc_hd__o21ai_1
X_5315_ _5546_/B vssd1 vssd1 vccd1 vccd1 _5514_/B sky130_fd_sc_hd__buf_2
X_5246_ _5246_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5177_ _5211_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5184_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _4470_/A _4470_/B _4470_/C vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__o21ai_2
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4059_ _4254_/A _4255_/A vssd1 vssd1 vccd1 vccd1 _4213_/D sky130_fd_sc_hd__and2_1
XFILLER_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6486__68 vssd1 vssd1 vccd1 vccd1 _6486__68/HI _6594_/A sky130_fd_sc_hd__conb_1
XFILLER_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3430_ _4886_/A _3430_/B _3430_/C vssd1 vssd1 vccd1 vccd1 _3449_/A sky130_fd_sc_hd__and3_1
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3361_ _5815_/A _4636_/A _6344_/Q vssd1 vssd1 vccd1 vccd1 _3364_/A sky130_fd_sc_hd__or3b_2
X_5100_ _5100_/A _5128_/B _5129_/A vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__and3_1
X_6080_ _6078_/X _6083_/B _6036_/A vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__a21bo_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5031_ _5031_/A _5045_/A vssd1 vssd1 vccd1 vccd1 _5045_/B sky130_fd_sc_hd__nand2_1
X_3292_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3297_/A sky130_fd_sc_hd__buf_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _5931_/X _5933_/B _5933_/C vssd1 vssd1 vccd1 vccd1 _5933_/X sky130_fd_sc_hd__and3b_1
X_5864_ _5846_/Y _5857_/X _5863_/X vssd1 vssd1 vccd1 vccd1 _6579_/A sky130_fd_sc_hd__o21a_1
X_4815_ _4820_/C _4815_/B vssd1 vssd1 vccd1 vccd1 _4816_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5795_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__buf_2
X_4746_ _3612_/A _4761_/B _4895_/D _4745_/X vssd1 vssd1 vccd1 vccd1 _4747_/C sky130_fd_sc_hd__a31o_1
XFILLER_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4677_ _4677_/A _4895_/D vssd1 vssd1 vccd1 vccd1 _4678_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6416_ _6423_/CLK _6416_/D vssd1 vssd1 vccd1 vccd1 _6416_/Q sky130_fd_sc_hd__dfxtp_1
X_3628_ _6327_/Q _6326_/Q _3628_/C _4694_/B vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__and4_1
X_6347_ _6426_/CLK _6347_/D vssd1 vssd1 vccd1 vccd1 _6347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3559_ _3565_/A _3565_/B vssd1 vssd1 vccd1 vccd1 _3563_/C sky130_fd_sc_hd__nand2_1
X_6278_ _6299_/A _6278_/B _6283_/C vssd1 vssd1 vccd1 vccd1 _6412_/D sky130_fd_sc_hd__nor3_1
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5229_ _5225_/A _5223_/X _5221_/X _5222_/X vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__o211a_1
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4600_ _5777_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4602_/A sky130_fd_sc_hd__xor2_1
X_5580_ _5384_/B _5580_/B vssd1 vssd1 vccd1 vccd1 _5580_/X sky130_fd_sc_hd__and2b_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4531_ _4523_/X _4522_/Y _4520_/Y vssd1 vssd1 vccd1 vccd1 _4531_/Y sky130_fd_sc_hd__a21oi_1
X_4462_ _4527_/A _4527_/B _4461_/X vssd1 vssd1 vccd1 vccd1 _4519_/B sky130_fd_sc_hd__a21o_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3413_ _3466_/A _3509_/B vssd1 vssd1 vccd1 vccd1 _3421_/B sky130_fd_sc_hd__nand2_1
X_6201_ _6376_/Q _6375_/Q _6378_/Q vssd1 vssd1 vccd1 vccd1 _6203_/B sky130_fd_sc_hd__or3_1
X_4393_ _5471_/C _4393_/B vssd1 vssd1 vccd1 vccd1 _4394_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3344_ _4272_/A vssd1 vssd1 vccd1 vccd1 _4104_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6132_ _6130_/X _6131_/X _6356_/Q _6100_/A vssd1 vssd1 vccd1 vccd1 _6132_/X sky130_fd_sc_hd__o211a_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3278_/A vssd1 vssd1 vccd1 vccd1 _3275_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6063_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6063_/Y sky130_fd_sc_hd__nand2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5014_ _5028_/A _5040_/B _5001_/B _5013_/X vssd1 vssd1 vccd1 vccd1 _5027_/B sky130_fd_sc_hd__a31o_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5916_ _5916_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5917_/B sky130_fd_sc_hd__or2_1
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5847_ _6416_/Q vssd1 vssd1 vccd1 vccd1 _5847_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5778_ _5778_/A _5778_/B vssd1 vssd1 vccd1 vccd1 _5779_/B sky130_fd_sc_hd__and2_1
X_4729_ _4728_/A _4812_/B _4728_/C vssd1 vssd1 vccd1 vccd1 _4730_/B sky130_fd_sc_hd__a21oi_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6456__38 vssd1 vssd1 vccd1 vccd1 _6456__38/HI _6561_/A sky130_fd_sc_hd__conb_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6470__52 vssd1 vssd1 vccd1 vccd1 _6470__52/HI _6575_/A sky130_fd_sc_hd__conb_1
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _4169_/C vssd1 vssd1 vccd1 vccd1 _4342_/B sky130_fd_sc_hd__clkbuf_2
X_5701_ _5702_/A _5702_/B vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__and2_1
X_3893_ _3893_/A _3893_/B vssd1 vssd1 vccd1 vccd1 _3917_/A sky130_fd_sc_hd__nor2_1
X_5632_ _5748_/A _5674_/A vssd1 vssd1 vccd1 vccd1 _5633_/B sky130_fd_sc_hd__xor2_1
X_5563_ _5706_/A _5698_/B vssd1 vssd1 vccd1 vccd1 _5699_/A sky130_fd_sc_hd__and2_1
XFILLER_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4514_ _4514_/A _4514_/B vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__and2_1
X_5494_ _5494_/A _5494_/B vssd1 vssd1 vccd1 vccd1 _5505_/A sky130_fd_sc_hd__xor2_1
XFILLER_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4445_ _4445_/A _4445_/B vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__nor2_1
X_4376_ _4377_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4380_/B sky130_fd_sc_hd__xor2_4
X_3327_ _3327_/A vssd1 vssd1 vccd1 vccd1 _3327_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6349_/Q _6115_/B vssd1 vssd1 vccd1 vccd1 _6116_/A sky130_fd_sc_hd__and2_1
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3260_/A vssd1 vssd1 vccd1 vccd1 _3258_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6338_/Q _6046_/B vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__or2_1
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4230_ _6323_/Q _5441_/A _4330_/B _4383_/C vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__and4_1
X_4161_ _4161_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4092_ _4072_/A _4072_/B _4072_/C vssd1 vssd1 vccd1 vccd1 _4113_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _5061_/B _5007_/A vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__nor2_1
X_3945_ _5006_/A _3958_/B _3959_/B _3944_/A vssd1 vssd1 vccd1 vccd1 _3947_/B sky130_fd_sc_hd__a31o_1
X_3876_ _5006_/A _4154_/B _3876_/C vssd1 vssd1 vccd1 vccd1 _3893_/A sky130_fd_sc_hd__and3_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5615_ _5615_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5615_/X sky130_fd_sc_hd__or2b_1
X_6595_ _6595_/A _3289_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5546_ _5546_/A _5546_/B vssd1 vssd1 vccd1 vccd1 _5547_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5477_ _5497_/A _5497_/B _5474_/A vssd1 vssd1 vccd1 vccd1 _5479_/B sky130_fd_sc_hd__o21ai_2
X_4428_ _5386_/A _4436_/B _5532_/B vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4359_ _4383_/A _4387_/B _4408_/B vssd1 vssd1 vccd1 vccd1 _4369_/B sky130_fd_sc_hd__and3_1
XFILLER_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _6401_/Q _6392_/Q vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__and2b_1
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6440__22 vssd1 vssd1 vccd1 vccd1 _6440__22/HI _6545_/A sky130_fd_sc_hd__conb_1
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3730_/A _3736_/A _3730_/C vssd1 vssd1 vccd1 vccd1 _3731_/C sky130_fd_sc_hd__nand3_1
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3661_ _3682_/A _3682_/B _3682_/C vssd1 vssd1 vccd1 vccd1 _3690_/A sky130_fd_sc_hd__a21oi_4
X_5400_ _5400_/A _5400_/B vssd1 vssd1 vccd1 vccd1 _5416_/B sky130_fd_sc_hd__xor2_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6380_ _6388_/CLK _6380_/D vssd1 vssd1 vccd1 vccd1 _6380_/Q sky130_fd_sc_hd__dfxtp_1
X_3592_ _4830_/B _4855_/A _3592_/C _3592_/D vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__nand4_4
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5331_ _5339_/B _5331_/B vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__xor2_4
XFILLER_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5262_ _5262_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__or2_1
X_4213_ _5407_/A _5387_/A _4213_/C _4213_/D vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__and4_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5193_ _5193_/A _5193_/B _5230_/A vssd1 vssd1 vccd1 vccd1 _5492_/C sky130_fd_sc_hd__or3b_4
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4144_ _4144_/A _4144_/B vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4075_ _4075_/A _4075_/B _4075_/C vssd1 vssd1 vccd1 vccd1 _4122_/A sky130_fd_sc_hd__and3_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4977_ _4977_/A _4977_/B vssd1 vssd1 vccd1 vccd1 _4995_/B sky130_fd_sc_hd__xnor2_4
X_3928_ _3928_/A _3928_/B vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__nor2_1
X_3859_ _6319_/Q vssd1 vssd1 vccd1 vccd1 _5487_/A sky130_fd_sc_hd__clkbuf_2
X_6578_ _6578_/A _3268_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5529_ _5570_/A _5570_/B vssd1 vssd1 vccd1 vccd1 _5529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4900_ _4900_/A _4900_/B vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__xnor2_1
X_5880_ _6419_/Q vssd1 vssd1 vccd1 vccd1 _6298_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4831_ _4831_/A _4831_/B _4842_/A vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__and3_1
X_4762_ _4762_/A _5997_/A _4755_/C vssd1 vssd1 vccd1 vccd1 _4805_/C sky130_fd_sc_hd__or3b_1
X_3713_ _3761_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__xor2_4
X_4693_ _4679_/A _4679_/B _4692_/X vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__o21ba_1
X_3644_ _3644_/A _3644_/B vssd1 vssd1 vccd1 vccd1 _3765_/B sky130_fd_sc_hd__xnor2_2
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3575_ _4697_/A _3589_/A _3534_/D _4802_/A vssd1 vssd1 vccd1 vccd1 _3576_/B sky130_fd_sc_hd__a22oi_1
X_6363_ _6396_/CLK _6363_/D vssd1 vssd1 vccd1 vccd1 _6363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5314_ _5486_/B vssd1 vssd1 vccd1 vccd1 _5546_/B sky130_fd_sc_hd__clkbuf_2
X_6294_ _6294_/A _6294_/B vssd1 vssd1 vccd1 vccd1 _6418_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _5245_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5176_ _5288_/B vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4127_ _4127_/A _4127_/B vssd1 vssd1 vccd1 vccd1 _4470_/C sky130_fd_sc_hd__nor2_1
XFILLER_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4058_ _4057_/A _4057_/B _3758_/X vssd1 vssd1 vccd1 vccd1 _4255_/A sky130_fd_sc_hd__o21bai_4
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6426_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3360_ _3409_/B vssd1 vssd1 vccd1 vccd1 _4636_/A sky130_fd_sc_hd__inv_2
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5030_ _5030_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__and2_1
X_3291_ _3291_/A vssd1 vssd1 vccd1 vccd1 _3291_/Y sky130_fd_sc_hd__inv_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5932_ _5761_/A _5765_/X _5829_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5933_/C sky130_fd_sc_hd__a31o_1
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5863_ _5847_/Y _5852_/X _5856_/Y _5858_/Y _6228_/A vssd1 vssd1 vccd1 vccd1 _5863_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _4814_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4815_/B sky130_fd_sc_hd__nand2_1
X_5794_ _5784_/A _5783_/Y _5792_/X _6405_/Q _5793_/X vssd1 vssd1 vccd1 vccd1 _5794_/X
+ sky130_fd_sc_hd__o221a_1
X_4745_ _4745_/A _4745_/B _4851_/A vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__and3_1
X_4676_ _4830_/D vssd1 vssd1 vccd1 vccd1 _4895_/D sky130_fd_sc_hd__clkbuf_2
X_6415_ _6423_/CLK _6415_/D vssd1 vssd1 vccd1 vccd1 _6415_/Q sky130_fd_sc_hd__dfxtp_1
X_3627_ _3627_/A _3627_/B vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__xor2_2
XFILLER_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3558_ _3558_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _3565_/B sky130_fd_sc_hd__xor2_1
X_6346_ _6361_/CLK _6346_/D vssd1 vssd1 vccd1 vccd1 _6346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3489_ _3489_/A _3489_/B vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__or2_1
X_6277_ _6412_/Q _6411_/Q _6410_/Q vssd1 vssd1 vccd1 vccd1 _6283_/C sky130_fd_sc_hd__and3_1
X_5228_ _5228_/A _5228_/B vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__nand2_4
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5159_ _5159_/A _5460_/B vssd1 vssd1 vccd1 vccd1 _5195_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4530_ _4523_/X _4520_/Y _4522_/Y _4528_/X _4529_/Y vssd1 vssd1 vccd1 vccd1 _4530_/X
+ sky130_fd_sc_hd__a32o_1
X_4461_ _4325_/B _4461_/B vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3412_ _3534_/D vssd1 vssd1 vccd1 vccd1 _3509_/B sky130_fd_sc_hd__clkbuf_2
X_6200_ _6376_/Q _6375_/Q _6378_/Q _6377_/Q vssd1 vssd1 vccd1 vccd1 _6200_/X sky130_fd_sc_hd__and4_1
XFILLER_98_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4392_ _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__xnor2_1
X_6131_ _6351_/Q _6352_/Q _6354_/Q _6353_/Q vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__or4_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _6323_/Q vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__clkbuf_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6062_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__or2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3278_/A vssd1 vssd1 vccd1 vccd1 _3274_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5013_ _5015_/A _5214_/B _5013_/C vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__and3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5915_ _5916_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__and2_1
X_5846_ _5838_/X _5841_/X _5845_/X vssd1 vssd1 vccd1 vccd1 _5846_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _5777_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _5778_/B sky130_fd_sc_hd__or2_1
X_4728_ _4728_/A _4728_/B _4728_/C vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__and3_1
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4659_ _4762_/A _4659_/B _4755_/C vssd1 vssd1 vccd1 vccd1 _4828_/A sky130_fd_sc_hd__and3b_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _6361_/CLK _6329_/D vssd1 vssd1 vccd1 vccd1 _6329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6523__105 vssd1 vssd1 vccd1 vccd1 _6523__105/HI _6631_/A sky130_fd_sc_hd__conb_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3961_/A _3961_/B vssd1 vssd1 vccd1 vccd1 _4169_/C sky130_fd_sc_hd__xor2_4
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5700_ _5700_/A vssd1 vssd1 vccd1 vccd1 _5702_/B sky130_fd_sc_hd__inv_2
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3892_ _5006_/A _4154_/B _3876_/C vssd1 vssd1 vccd1 vccd1 _3893_/B sky130_fd_sc_hd__a21oi_1
X_5631_ _5681_/A _5803_/A vssd1 vssd1 vccd1 vccd1 _5633_/A sky130_fd_sc_hd__nor2_1
X_5562_ _5692_/A _5562_/B vssd1 vssd1 vccd1 vccd1 _5698_/B sky130_fd_sc_hd__nor2_1
X_4513_ _5777_/B _4513_/B vssd1 vssd1 vccd1 vccd1 _4514_/B sky130_fd_sc_hd__and2_1
X_5493_ _5495_/B _5493_/B vssd1 vssd1 vccd1 vccd1 _5509_/A sky130_fd_sc_hd__and2b_1
X_4444_ _4575_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__or2_1
X_4375_ _5471_/C _4372_/A _4393_/B _4381_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4377_/B
+ sky130_fd_sc_hd__a32o_2
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3326_ _3327_/A vssd1 vssd1 vccd1 vccd1 _3326_/Y sky130_fd_sc_hd__inv_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6114_/A vssd1 vssd1 vccd1 vccd1 _6349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6338_/Q _6059_/A vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__nand2_1
X_3257_ _3260_/A vssd1 vssd1 vccd1 vccd1 _3257_/Y sky130_fd_sc_hd__inv_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5829_ _5829_/A vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6516__98 vssd1 vssd1 vccd1 vccd1 _6516__98/HI _6624_/A sky130_fd_sc_hd__conb_1
XFILLER_77_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4160_ _4160_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _4160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ _4089_/A _4087_/X _4079_/C _4086_/Y vssd1 vssd1 vccd1 vccd1 _4470_/B sky130_fd_sc_hd__o211a_1
XFILLER_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4993_ _5060_/A _5096_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ _3944_/A _3944_/B vssd1 vssd1 vccd1 vccd1 _3959_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3875_ _3875_/A _3898_/A vssd1 vssd1 vccd1 vccd1 _3876_/C sky130_fd_sc_hd__xor2_1
X_5614_ _5602_/A _5602_/B _5605_/B vssd1 vssd1 vccd1 vccd1 _5614_/X sky130_fd_sc_hd__a21o_1
X_6594_ _6594_/A _3288_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5545_ _5545_/A _5545_/B _5545_/C vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__and3_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5476_ _5476_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5497_/B sky130_fd_sc_hd__xnor2_2
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4427_ _5545_/C vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4358_ _6319_/Q _4383_/C vssd1 vssd1 vccd1 vccd1 _4408_/B sky130_fd_sc_hd__and2_1
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4289_ _4262_/A _4262_/B _4288_/Y vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__o21ba_1
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3309_/Y sky130_fd_sc_hd__inv_2
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6028_ _6334_/Q _6355_/Q vssd1 vssd1 vccd1 vccd1 _6028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6529__111 vssd1 vssd1 vccd1 vccd1 _6529__111/HI _6637_/A sky130_fd_sc_hd__conb_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3660_ _3660_/A _3660_/B vssd1 vssd1 vccd1 vccd1 _3682_/C sky130_fd_sc_hd__or2_1
X_3591_ _3591_/A _3591_/B vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__xnor2_2
X_5330_ _5330_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _5331_/B sky130_fd_sc_hd__xnor2_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5261_ _5267_/B _5261_/B vssd1 vssd1 vccd1 vccd1 _5272_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4212_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__nand2_1
X_5192_ _5192_/A _5192_/B vssd1 vssd1 vccd1 vccd1 _5226_/A sky130_fd_sc_hd__xor2_1
XFILLER_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4143_ _4143_/A _4143_/B vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4074_ _4075_/A _4075_/B _4075_/C vssd1 vssd1 vccd1 vccd1 _4074_/Y sky130_fd_sc_hd__nand3_1
XFILLER_83_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _4974_/A _4974_/B _4939_/Y vssd1 vssd1 vccd1 vccd1 _4977_/A sky130_fd_sc_hd__o21a_1
XFILLER_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3927_ _3927_/A _3927_/B vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__and2_1
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3858_ _5015_/A _3858_/B vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__nand2_1
X_3789_ _3931_/A vssd1 vssd1 vccd1 vccd1 _3818_/B sky130_fd_sc_hd__buf_2
X_6577_ _6577_/A _3266_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
X_5528_ _5530_/A _5530_/B _5527_/X vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__o21a_1
XFILLER_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5459_ _5476_/A _5457_/X _5458_/X vssd1 vssd1 vccd1 vccd1 _5460_/C sky130_fd_sc_hd__a21o_1
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6500__82 vssd1 vssd1 vccd1 vccd1 _6500__82/HI _6608_/A sky130_fd_sc_hd__conb_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4830_ _4830_/A _4830_/B _4830_/C _4830_/D vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__nand4_4
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _4745_/X _4761_/B vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__and2b_1
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3712_ _3712_/A _3759_/A vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__nand2_2
X_4692_ _4711_/A _4891_/D _4692_/C vssd1 vssd1 vccd1 vccd1 _4692_/X sky130_fd_sc_hd__and3_1
X_3643_ _3767_/A _3767_/B vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__xor2_4
X_6362_ _6396_/CLK _6362_/D vssd1 vssd1 vccd1 vccd1 _6362_/Q sky130_fd_sc_hd__dfxtp_1
X_3574_ _3716_/C vssd1 vssd1 vccd1 vccd1 _3589_/A sky130_fd_sc_hd__clkbuf_2
X_5313_ _5313_/A _5313_/B vssd1 vssd1 vccd1 vccd1 _5486_/B sky130_fd_sc_hd__xnor2_1
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6293_ _6417_/Q _6290_/B _6292_/Y vssd1 vssd1 vccd1 vccd1 _6417_/D sky130_fd_sc_hd__o21a_1
XFILLER_115_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5244_ _5244_/A _5244_/B _5274_/A vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__nor3_1
X_5175_ _5175_/A _5175_/B _5174_/Y vssd1 vssd1 vccd1 vccd1 _5219_/B sky130_fd_sc_hd__or3b_1
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4118_/C _4121_/B _4127_/A _4125_/X vssd1 vssd1 vccd1 vccd1 _4127_/B sky130_fd_sc_hd__a211oi_4
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ _4057_/A _4057_/B _3758_/X vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__or3b_2
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4959_ _5313_/A _4959_/B vssd1 vssd1 vccd1 vccd1 _4960_/B sky130_fd_sc_hd__or2_1
XFILLER_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6629_ _6629_/A _3327_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3290_ _3291_/A vssd1 vssd1 vccd1 vccd1 _3290_/Y sky130_fd_sc_hd__inv_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6477__59 vssd1 vssd1 vccd1 vccd1 _6477__59/HI _6585_/A sky130_fd_sc_hd__conb_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5931_ _5761_/A _5927_/A _5944_/A vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5862_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6228_/A sky130_fd_sc_hd__buf_2
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4813_ _4813_/A _4813_/B vssd1 vssd1 vccd1 vccd1 _4820_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5793_ _6404_/Q _5793_/B vssd1 vssd1 vccd1 vccd1 _5793_/X sky130_fd_sc_hd__or2_1
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4744_ _6333_/Q _4805_/B _4830_/C _3647_/A vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__a22o_1
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4675_ _4690_/A vssd1 vssd1 vccd1 vccd1 _4830_/D sky130_fd_sc_hd__clkbuf_2
X_3626_ _3626_/A _3626_/B vssd1 vssd1 vccd1 vccd1 _3635_/A sky130_fd_sc_hd__xnor2_2
X_6414_ _6426_/CLK _6414_/D vssd1 vssd1 vccd1 vccd1 _6414_/Q sky130_fd_sc_hd__dfxtp_1
X_3557_ _3529_/B _3576_/A _3529_/A vssd1 vssd1 vccd1 vccd1 _3565_/A sky130_fd_sc_hd__o21bai_1
X_6345_ _6345_/CLK _6345_/D vssd1 vssd1 vccd1 vccd1 _6345_/Q sky130_fd_sc_hd__dfxtp_1
X_6276_ _5828_/X _6273_/A _6412_/Q vssd1 vssd1 vccd1 vccd1 _6278_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5227_ _5227_/A _5226_/A vssd1 vssd1 vccd1 vccd1 _5228_/B sky130_fd_sc_hd__or2b_1
X_3488_ _4697_/B _3406_/B _3430_/B _4802_/A vssd1 vssd1 vccd1 vccd1 _3489_/B sky130_fd_sc_hd__a22oi_1
X_5158_ _5322_/B vssd1 vssd1 vccd1 vccd1 _5460_/B sky130_fd_sc_hd__buf_2
X_4109_ _4109_/A _4109_/B _4109_/C vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__and3_1
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5089_ _5090_/B _5090_/C _5090_/A vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__o21a_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491__73 vssd1 vssd1 vccd1 vccd1 _6491__73/HI _6599_/A sky130_fd_sc_hd__conb_1
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _4572_/A _4572_/B _4459_/X vssd1 vssd1 vccd1 vccd1 _4527_/B sky130_fd_sc_hd__a21o_2
XFILLER_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4391_ _5492_/A _4391_/B _4391_/C vssd1 vssd1 vccd1 vccd1 _4397_/B sky130_fd_sc_hd__and3_1
X_3411_ _3650_/B vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__clkbuf_2
X_3342_ _3342_/A vssd1 vssd1 vccd1 vccd1 _3342_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6130_ _6347_/Q _6348_/Q _6349_/Q _6350_/Q vssd1 vssd1 vccd1 vccd1 _6130_/X sky130_fd_sc_hd__or4_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3279_/A vssd1 vssd1 vccd1 vccd1 _3278_/A sky130_fd_sc_hd__buf_12
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6052_/X _6056_/B _6054_/B vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__o21a_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5012_ _5113_/B vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__buf_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5914_ _5902_/X _5904_/X _5905_/X _5903_/Y vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__o22a_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5845_ _6414_/Q _5840_/Y _5844_/Y _6415_/Q vssd1 vssd1 vccd1 vccd1 _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5776_ _5776_/A _5776_/B vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__or2_1
X_4727_ _4697_/A _4854_/B _4769_/B _4697_/B vssd1 vssd1 vccd1 vccd1 _4728_/C sky130_fd_sc_hd__a22o_1
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4658_ _3356_/A _6345_/Q _6337_/Q _6336_/Q vssd1 vssd1 vccd1 vccd1 _4755_/C sky130_fd_sc_hd__a211o_1
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3609_ _6329_/Q vssd1 vssd1 vccd1 vccd1 _4755_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4589_ _4565_/A _4565_/B _4587_/X _4588_/Y vssd1 vssd1 vccd1 vccd1 _4589_/X sky130_fd_sc_hd__a22o_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6328_ _6361_/CLK _6328_/D vssd1 vssd1 vccd1 vccd1 _6328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6405_/Q _6262_/C vssd1 vssd1 vccd1 vccd1 _6260_/B sky130_fd_sc_hd__and2_1
XFILLER_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6447__29 vssd1 vssd1 vccd1 vccd1 _6447__29/HI _6552_/A sky130_fd_sc_hd__conb_1
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3960_ _3960_/A _4302_/B vssd1 vssd1 vccd1 vccd1 _3960_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ _3891_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__xor2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5630_ _5630_/A _5630_/B vssd1 vssd1 vccd1 vccd1 _5681_/A sky130_fd_sc_hd__xnor2_4
XFILLER_31_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5561_ _5428_/A _5555_/D _5547_/B _5554_/Y vssd1 vssd1 vccd1 vccd1 _5562_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5492_ _5492_/A _5492_/B _5492_/C vssd1 vssd1 vccd1 vccd1 _5493_/B sky130_fd_sc_hd__and3_1
X_4512_ _4618_/A _4512_/B vssd1 vssd1 vccd1 vccd1 _4513_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4443_ _4443_/A _4443_/B vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__or2_1
X_4374_ _4374_/A _4374_/B vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__xnor2_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3327_/A vssd1 vssd1 vccd1 vccd1 _3325_/Y sky130_fd_sc_hd__inv_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6348_/Q _6234_/A vssd1 vssd1 vccd1 vccd1 _6114_/A sky130_fd_sc_hd__and2_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3256_ _3260_/A vssd1 vssd1 vccd1 vccd1 _3256_/Y sky130_fd_sc_hd__inv_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6046_/B vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461__43 vssd1 vssd1 vccd1 vccd1 _6461__43/HI _6566_/A sky130_fd_sc_hd__conb_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5828_ _6411_/Q vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5759_ _5759_/A _5789_/B vssd1 vssd1 vccd1 vccd1 _5759_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4090_ _4472_/A _4472_/B _4472_/C vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4992_ _5202_/B vssd1 vssd1 vccd1 vccd1 _5096_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ _3943_/A _3966_/A vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__and2_1
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3874_ _5433_/A _3958_/B vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__nand2_1
X_5613_ _5613_/A _5613_/B vssd1 vssd1 vccd1 vccd1 _5796_/A sky130_fd_sc_hd__xnor2_4
X_6593_ _6593_/A _3287_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
X_5544_ _5544_/A _5544_/B vssd1 vssd1 vccd1 vccd1 _5556_/A sky130_fd_sc_hd__xor2_1
X_5475_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5476_/B sky130_fd_sc_hd__xor2_1
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4426_ _4431_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__or2_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4357_ _5424_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__nand2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4288_/A _4288_/B vssd1 vssd1 vccd1 vccd1 _4288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3308_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__inv_2
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3241_/A vssd1 vssd1 vccd1 vccd1 _3239_/Y sky130_fd_sc_hd__inv_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6334_/Q _6355_/Q vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__and2_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3590_ _6010_/A _3589_/Y _3573_/B vssd1 vssd1 vccd1 vccd1 _3626_/A sky130_fd_sc_hd__o21a_1
XFILLER_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5260_ _5296_/A _5350_/B _5259_/C vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__a21o_1
X_4211_ _5387_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4211_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5191_ _5191_/A _5191_/B _5191_/C vssd1 vssd1 vccd1 vccd1 _5647_/A sky130_fd_sc_hd__and3_2
X_4142_ _5350_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4143_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4073_ _4071_/A _4071_/B _4113_/A vssd1 vssd1 vccd1 vccd1 _4075_/C sky130_fd_sc_hd__a21o_1
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6431__13 vssd1 vssd1 vccd1 vccd1 _6431__13/HI _6536_/A sky130_fd_sc_hd__conb_1
X_4975_ _4987_/A _4987_/B _4975_/C vssd1 vssd1 vccd1 vccd1 _4995_/A sky130_fd_sc_hd__or3_4
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3926_ _3927_/A _3927_/B vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__nor2_1
X_3857_ _3857_/A _3857_/B vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__or2_1
X_3788_ _3788_/A _3788_/B vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__xnor2_4
X_6576_ _6576_/A _3265_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_5527_ _5527_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5527_/X sky130_fd_sc_hd__or2b_1
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5458_ _5458_/A _5458_/B _5475_/B vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__and3_1
X_5389_ _5425_/A _5460_/B vssd1 vssd1 vccd1 vccd1 _5401_/B sky130_fd_sc_hd__nand2_1
X_4409_ _4409_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__nor2_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4760_ _4888_/A _4758_/B _4770_/A _4758_/D vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3711_ _3712_/A _3711_/B _3711_/C vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__nand3_2
X_4691_ _4850_/B vssd1 vssd1 vccd1 vccd1 _4891_/D sky130_fd_sc_hd__clkbuf_2
X_3642_ _3642_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3767_/B sky130_fd_sc_hd__and2_2
X_6361_ _6361_/CLK _6361_/D vssd1 vssd1 vccd1 vccd1 _6361_/Q sky130_fd_sc_hd__dfxtp_1
X_3573_ _3573_/A _3573_/B vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__nand2_1
X_5312_ _5369_/A _5368_/A _4959_/B vssd1 vssd1 vccd1 vccd1 _5313_/B sky130_fd_sc_hd__a21bo_1
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6292_ _6417_/Q _6290_/B _6007_/X vssd1 vssd1 vccd1 vccd1 _6292_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5243_ _5244_/B _5274_/A _5244_/A vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__o21a_1
X_5174_ _5174_/A _5174_/B vssd1 vssd1 vccd1 vccd1 _5174_/Y sky130_fd_sc_hd__xnor2_1
X_4125_ _4122_/Y _4123_/X _4121_/A _4121_/Y vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__o211a_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4056_ _3759_/A _3759_/B _3759_/C vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__a21oi_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4958_ _5369_/A _5368_/B vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__or2b_1
X_3909_ _5458_/A vssd1 vssd1 vccd1 vccd1 _5350_/A sky130_fd_sc_hd__clkbuf_2
X_4889_ _4886_/Y _4888_/Y _4875_/B vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__a21oi_1
X_6628_ _6628_/A _3326_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6559_ _6559_/A _3245_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5930_ _5930_/A vssd1 vssd1 vccd1 vccd1 _6318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5861_ _6025_/B vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4812_ _4956_/A _4812_/B vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5792_ _5785_/X _5746_/X _5791_/X _5743_/A vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4743_ _4745_/B vssd1 vssd1 vccd1 vccd1 _4830_/C sky130_fd_sc_hd__clkbuf_2
X_6413_ _6426_/CLK _6413_/D vssd1 vssd1 vccd1 vccd1 _6413_/Q sky130_fd_sc_hd__dfxtp_1
X_4674_ _4755_/C _3607_/A _4648_/B vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__a21boi_1
X_3625_ _3625_/A _3625_/B vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__or2_1
X_3556_ _3558_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__or2_1
X_6344_ _6361_/CLK _6344_/D vssd1 vssd1 vccd1 vccd1 _6344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6275_ _5828_/X _6273_/A _6274_/Y vssd1 vssd1 vccd1 vccd1 _6411_/D sky130_fd_sc_hd__a21oi_1
X_5226_ _5226_/A _5227_/A vssd1 vssd1 vccd1 vccd1 _5228_/A sky130_fd_sc_hd__or2b_2
X_3487_ _4850_/A vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5157_ _5492_/B _5157_/B vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__xnor2_1
X_4108_ _4110_/B _4108_/B vssd1 vssd1 vccd1 vccd1 _4109_/C sky130_fd_sc_hd__nor2_1
X_5088_ _5088_/A _5088_/B vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__and2_1
X_4039_ _4022_/B _4037_/Y _5121_/A _4079_/B vssd1 vssd1 vccd1 vccd1 _4047_/A sky130_fd_sc_hd__o211ai_2
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4390_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__xnor2_1
X_3410_ _6342_/Q _3472_/B vssd1 vssd1 vccd1 vccd1 _3650_/B sky130_fd_sc_hd__or2_2
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3341_ _3342_/A vssd1 vssd1 vccd1 vccd1 _3341_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3272_ _3272_/A vssd1 vssd1 vccd1 vccd1 _3272_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6060_ _6060_/A _6074_/B vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__xor2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5011_ _5075_/A _5074_/B _5074_/A vssd1 vssd1 vccd1 vccd1 _5022_/B sky130_fd_sc_hd__o21ba_1
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5913_ _5918_/A _5909_/X _5912_/Y vssd1 vssd1 vccd1 vccd1 _6316_/D sky130_fd_sc_hd__a21oi_1
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5844_ _5945_/A _5825_/X _5843_/X _5807_/X vssd1 vssd1 vccd1 vccd1 _5844_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5775_ _5775_/A _5775_/B vssd1 vssd1 vccd1 vccd1 _5775_/Y sky130_fd_sc_hd__nor2_1
X_4726_ _4834_/B vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4657_ _3356_/A _3359_/A _6337_/Q _6336_/Q vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__a22o_1
X_3608_ _3646_/A _3646_/C _3699_/D vssd1 vssd1 vccd1 vccd1 _3608_/Y sky130_fd_sc_hd__nand3_1
X_4588_ _4588_/A _4588_/B vssd1 vssd1 vccd1 vccd1 _4588_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6327_ _6345_/CLK _6327_/D vssd1 vssd1 vccd1 vccd1 _6327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3539_ _4850_/A _3538_/X _3547_/A vssd1 vssd1 vccd1 vccd1 _3591_/A sky130_fd_sc_hd__a21boi_4
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6258_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6280_/A sky130_fd_sc_hd__buf_2
XFILLER_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5209_ _5210_/A _5210_/B vssd1 vssd1 vccd1 vccd1 _5209_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6189_ _6189_/A vssd1 vssd1 vccd1 vccd1 _6378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3890_ _3890_/A _3890_/B vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__and2_1
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5560_ _5560_/A _5560_/B _5560_/C vssd1 vssd1 vccd1 vccd1 _5706_/A sky130_fd_sc_hd__and3_1
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4511_ _4540_/A _5750_/A vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__and2b_1
X_5491_ _5488_/A _5511_/A _5490_/X vssd1 vssd1 vccd1 vccd1 _5495_/B sky130_fd_sc_hd__o21a_1
X_4442_ _4441_/B _4441_/C _4441_/A vssd1 vssd1 vccd1 vccd1 _4443_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4373_ _4373_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4374_/A sky130_fd_sc_hd__nand2_2
X_3324_ _3327_/A vssd1 vssd1 vccd1 vccd1 _3324_/Y sky130_fd_sc_hd__inv_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6126_/B vssd1 vssd1 vccd1 vccd1 _6234_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3255_ _3279_/A vssd1 vssd1 vccd1 vccd1 _3260_/A sky130_fd_sc_hd__buf_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6038_/A _6036_/X _6042_/Y _6015_/X vssd1 vssd1 vccd1 vccd1 _6337_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5827_ _5785_/X _5825_/X _5826_/Y _5743_/X vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__o2bb2a_1
X_5758_ _5758_/A _5767_/A vssd1 vssd1 vccd1 vccd1 _5758_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709_ _4749_/B vssd1 vssd1 vccd1 vccd1 _4834_/B sky130_fd_sc_hd__clkbuf_2
X_5689_ _5937_/A _5691_/B _5688_/Y vssd1 vssd1 vccd1 vccd1 _5723_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6507__89 vssd1 vssd1 vccd1 vccd1 _6507__89/HI _6615_/A sky130_fd_sc_hd__conb_1
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4991_ _4995_/A _4991_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__nand2_2
X_3942_ _3943_/A _3966_/A vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__nor2_1
X_3873_ _4221_/B vssd1 vssd1 vccd1 vccd1 _3958_/B sky130_fd_sc_hd__buf_2
XFILLER_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6592_ _6592_/A _3284_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_5612_ _5615_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5748_/A sky130_fd_sc_hd__xor2_4
X_5543_ _5543_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5565_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5474_ _5474_/A _5474_/B vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__nand2_1
X_4425_ _5546_/A _4406_/B _4188_/X _5514_/A vssd1 vssd1 vccd1 vccd1 _4426_/B sky130_fd_sc_hd__a22oi_1
X_4356_ _4356_/A vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__inv_2
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3307_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4287_ _4290_/B _4290_/A vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__and2b_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3238_ _3241_/A vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A vssd1 vssd1 vccd1 vccd1 _6335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4210_ _5456_/A vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__clkbuf_2
X_5190_ _5192_/B _5192_/A vssd1 vssd1 vccd1 vccd1 _5191_/C sky130_fd_sc_hd__or2b_1
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4141_ _4141_/A _4141_/B vssd1 vssd1 vccd1 vccd1 _4143_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _4072_/A _4072_/B _4072_/C vssd1 vssd1 vccd1 vccd1 _4113_/A sky130_fd_sc_hd__and3_1
XFILLER_95_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4974_ _4974_/A _4974_/B vssd1 vssd1 vccd1 vccd1 _4975_/C sky130_fd_sc_hd__xnor2_1
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3925_ _3925_/A _3925_/B vssd1 vssd1 vccd1 vccd1 _3927_/B sky130_fd_sc_hd__xnor2_1
X_3856_ _3856_/A _3856_/B vssd1 vssd1 vccd1 vccd1 _3857_/B sky130_fd_sc_hd__nor2_1
X_3787_ _3787_/A _3483_/X vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__or2b_2
X_6575_ _6575_/A _3264_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
X_5526_ _5527_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5530_/B sky130_fd_sc_hd__xor2_2
X_5457_ _5475_/A _5475_/B vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__or2_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4408_ _5545_/C _4408_/B _4424_/C vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__and3_1
X_5388_ _5390_/A _5390_/B vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__xnor2_2
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4339_ _4335_/A _4335_/B _4333_/B vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__a21o_2
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6009_ _4629_/A _6006_/X _6008_/Y vssd1 vssd1 vccd1 vccd1 _6331_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3710_ _3707_/A _3707_/B _3730_/A vssd1 vssd1 vccd1 vccd1 _3711_/C sky130_fd_sc_hd__a21o_1
X_4690_ _4690_/A vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__clkbuf_2
X_3641_ _3644_/A _3644_/B vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__or2b_1
X_3572_ _3525_/A _3716_/C _3589_/B vssd1 vssd1 vccd1 vccd1 _3573_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6360_ _6361_/CLK _6360_/D vssd1 vssd1 vccd1 vccd1 _6360_/Q sky130_fd_sc_hd__dfxtp_1
X_5311_ _5311_/A _5311_/B vssd1 vssd1 vccd1 vccd1 _5326_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6291_ _6416_/Q _6287_/B _6290_/Y vssd1 vssd1 vccd1 vccd1 _6416_/D sky130_fd_sc_hd__o21a_1
X_5242_ _5242_/A _5242_/B vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5173_ _5208_/A _5208_/B vssd1 vssd1 vccd1 vccd1 _5175_/B sky130_fd_sc_hd__and2_1
X_4124_ _4121_/A _4121_/Y _4122_/Y _4123_/X vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__a211oi_4
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4055_ _4055_/A _4055_/B vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4957_ _4957_/A _4957_/B _4957_/C vssd1 vssd1 vccd1 vccd1 _5368_/B sky130_fd_sc_hd__and3_1
X_3908_ _5386_/A vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__buf_2
X_4888_ _4888_/A _4956_/B vssd1 vssd1 vccd1 vccd1 _4888_/Y sky130_fd_sc_hd__nand2_1
X_6519__101 vssd1 vssd1 vccd1 vccd1 _6519__101/HI _6627_/A sky130_fd_sc_hd__conb_1
XFILLER_32_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3839_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5851_/A sky130_fd_sc_hd__clkbuf_4
X_6627_ _6627_/A _3325_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6558_ _6558_/A _3244_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5509_ _5509_/A _5509_/B vssd1 vssd1 vccd1 vccd1 _5570_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5860_ _6126_/B vssd1 vssd1 vccd1 vccd1 _6025_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4811_ _4811_/A _4811_/B vssd1 vssd1 vccd1 vccd1 _4826_/A sky130_fd_sc_hd__xnor2_2
X_5791_ _4639_/A _5788_/Y _5790_/Y _5751_/Y vssd1 vssd1 vccd1 vccd1 _5791_/X sky130_fd_sc_hd__o2bb2a_1
X_4742_ _3612_/A _4873_/B _4668_/A _4667_/D vssd1 vssd1 vccd1 vccd1 _4747_/B sky130_fd_sc_hd__a22o_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4672_/X _4673_/B _4751_/C vssd1 vssd1 vccd1 vccd1 _4692_/C sky130_fd_sc_hd__and3b_1
X_3624_ _3624_/A _3651_/A vssd1 vssd1 vccd1 vccd1 _3625_/B sky130_fd_sc_hd__nor2_1
X_6412_ _6426_/CLK _6412_/D vssd1 vssd1 vccd1 vccd1 _6412_/Q sky130_fd_sc_hd__dfxtp_1
X_3555_ _3585_/A _3585_/B _3554_/A vssd1 vssd1 vccd1 vccd1 _3558_/B sky130_fd_sc_hd__o21a_1
X_6343_ _6345_/CLK _6343_/D vssd1 vssd1 vccd1 vccd1 _6343_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6274_ _5828_/X _6273_/A _5911_/X vssd1 vssd1 vccd1 vccd1 _6274_/Y sky130_fd_sc_hd__o21ai_1
X_3486_ _6328_/Q vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__buf_2
X_5225_ _5225_/A _5225_/B vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__or2_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5156_ _5234_/A vssd1 vssd1 vccd1 vccd1 _5492_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4107_ _5237_/A _4212_/B _4412_/B _4104_/A vssd1 vssd1 vccd1 vccd1 _4108_/B sky130_fd_sc_hd__a22oi_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5087_ _5087_/A _5087_/B _5087_/C vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__or3_1
X_4038_ _5246_/A vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__buf_2
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _5985_/A _5982_/A _5988_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _6328_/D sky130_fd_sc_hd__o211a_1
XFILLER_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6482__64 vssd1 vssd1 vccd1 vccd1 _6482__64/HI _6590_/A sky130_fd_sc_hd__conb_1
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3340_ _3342_/A vssd1 vssd1 vccd1 vccd1 _3340_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6401_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5010_ _5009_/A _5009_/B _5009_/C vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__o21a_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3272_/A vssd1 vssd1 vccd1 vccd1 _3271_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5912_ _5918_/A _5954_/A _5911_/X vssd1 vssd1 vccd1 vccd1 _5912_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5843_ _5818_/X _5805_/X _5820_/X _5804_/X vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5774_ _5774_/A _5774_/B _5774_/C vssd1 vssd1 vccd1 vccd1 _5775_/B sky130_fd_sc_hd__and3_1
X_4725_ _4715_/A _4715_/B _4724_/X vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__o21a_1
XFILLER_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4656_ _4682_/A _4812_/B _4683_/B _4655_/Y vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__a31o_1
X_4587_ _4588_/A _4588_/B _4563_/Y _4586_/X vssd1 vssd1 vccd1 vccd1 _4587_/X sky130_fd_sc_hd__a2bb2o_1
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _3699_/D sky130_fd_sc_hd__clkbuf_2
X_6326_ _6345_/CLK _6326_/D vssd1 vssd1 vccd1 vccd1 _6326_/Q sky130_fd_sc_hd__dfxtp_1
X_3538_ _6326_/Q _4694_/B _3538_/C vssd1 vssd1 vccd1 vccd1 _3538_/X sky130_fd_sc_hd__and3_1
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3469_ _3469_/A _3469_/B _3469_/C vssd1 vssd1 vccd1 vccd1 _3470_/B sky130_fd_sc_hd__and3_1
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6294_/B _6257_/B _6262_/C vssd1 vssd1 vccd1 vccd1 _6404_/D sky130_fd_sc_hd__nor3_1
XFILLER_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5208_/A _5208_/B vssd1 vssd1 vccd1 vccd1 _5210_/B sky130_fd_sc_hd__xor2_2
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6188_ _6377_/Q _6194_/B vssd1 vssd1 vccd1 vccd1 _6189_/A sky130_fd_sc_hd__and2_1
XFILLER_97_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5139_ _5144_/A _5144_/B vssd1 vssd1 vccd1 vccd1 _5140_/B sky130_fd_sc_hd__xor2_1
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _4510_/A _4510_/B vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__xnor2_4
X_5490_ _5498_/A _5498_/B vssd1 vssd1 vccd1 vccd1 _5490_/X sky130_fd_sc_hd__or2_1
X_4441_ _4441_/A _4441_/B _4441_/C vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__and3_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4372_ _4372_/A _4394_/A vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__xor2_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6111_/A vssd1 vssd1 vccd1 vccd1 _6348_/D sky130_fd_sc_hd__clkbuf_1
X_3323_ _3327_/A vssd1 vssd1 vccd1 vccd1 _3323_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ input1/X vssd1 vssd1 vccd1 vccd1 _3279_/A sky130_fd_sc_hd__clkbuf_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6039_/X _6040_/Y _6099_/A vssd1 vssd1 vccd1 vccd1 _6042_/Y sky130_fd_sc_hd__o21ai_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5826_ _3364_/A _5790_/Y _5820_/X _5788_/Y vssd1 vssd1 vccd1 vccd1 _5826_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5757_ _5766_/B _5775_/A _5766_/A vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__o21ai_2
X_4708_ _4700_/A _4699_/B _4699_/A vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__o21ba_1
X_5688_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5688_/Y sky130_fd_sc_hd__nor2_1
X_4639_ _4639_/A vssd1 vssd1 vccd1 vccd1 _5742_/A sky130_fd_sc_hd__inv_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6309_ _6424_/Q _6423_/Q _6309_/C vssd1 vssd1 vccd1 vccd1 _6310_/B sky130_fd_sc_hd__and3_1
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6452__34 vssd1 vssd1 vccd1 vccd1 _6452__34/HI _6557_/A sky130_fd_sc_hd__conb_1
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4990_ _4987_/A _4987_/B _4975_/C vssd1 vssd1 vccd1 vccd1 _4991_/B sky130_fd_sc_hd__o21ai_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _4014_/A _4302_/B vssd1 vssd1 vccd1 vccd1 _3966_/A sky130_fd_sc_hd__nand2_1
X_3872_ _4068_/B vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6591_ _6591_/A _3283_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
X_5611_ _5613_/A _5613_/B _5600_/A _5610_/X vssd1 vssd1 vccd1 vccd1 _5612_/B sky130_fd_sc_hd__a31o_2
X_5542_ _5568_/A _5568_/B vssd1 vssd1 vccd1 vccd1 _5673_/A sky130_fd_sc_hd__xor2_2
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5473_ _5473_/A _5500_/A vssd1 vssd1 vccd1 vccd1 _5474_/B sky130_fd_sc_hd__or2_1
X_4424_ _5546_/A _4424_/B _4424_/C vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__and3_1
XFILLER_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4355_ _6319_/Q _4330_/B _4383_/C _4383_/A vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__a22o_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4286_ _4286_/A _4286_/B vssd1 vssd1 vccd1 vccd1 _4290_/A sky130_fd_sc_hd__xor2_1
XFILLER_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3241_/A vssd1 vssd1 vccd1 vccd1 _3237_/Y sky130_fd_sc_hd__inv_2
X_6025_ _6383_/Q _6025_/B vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__and2_1
XFILLER_67_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5809_ _6406_/Q _5800_/X _5808_/Y _6407_/Q vssd1 vssd1 vccd1 vccd1 _5809_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4140_ _5317_/A _4140_/B _4140_/C vssd1 vssd1 vccd1 vccd1 _4141_/B sky130_fd_sc_hd__and3_1
X_4071_ _4071_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4072_/C sky130_fd_sc_hd__xor2_1
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4973_ _4973_/A _4973_/B vssd1 vssd1 vccd1 vccd1 _4987_/B sky130_fd_sc_hd__xor2_2
X_3924_ _4476_/A _4476_/B vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3855_ _3855_/A _3855_/B vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__nand2_1
X_3786_ _5060_/A vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6574_ _6574_/A _3263_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_5525_ _5531_/A _5531_/B _5524_/Y vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__a21o_1
X_5456_ _5456_/A _5546_/B vssd1 vssd1 vccd1 vccd1 _5475_/B sky130_fd_sc_hd__and2_1
X_4407_ _5545_/C _4408_/B _4424_/C vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__a21oi_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5387_ _5387_/A _5455_/B _5455_/C vssd1 vssd1 vccd1 vccd1 _5390_/B sky130_fd_sc_hd__and3_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4338_/A _4338_/B vssd1 vssd1 vccd1 vccd1 _4368_/B sky130_fd_sc_hd__or2_2
XFILLER_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4269_ _6322_/Q vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__inv_4
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6008_ _4629_/A _6006_/X _6007_/X vssd1 vssd1 vccd1 vccd1 _6008_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3640_/A _3640_/B vssd1 vssd1 vccd1 vccd1 _3644_/B sky130_fd_sc_hd__xnor2_1
X_3571_ _3612_/A _3570_/X _3573_/A vssd1 vssd1 vccd1 vccd1 _3589_/B sky130_fd_sc_hd__a21bo_1
X_5310_ _5310_/A _5310_/B vssd1 vssd1 vccd1 vccd1 _5583_/A sky130_fd_sc_hd__xnor2_4
X_6290_ _6304_/A _6290_/B vssd1 vssd1 vccd1 vccd1 _6290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5241_ _5154_/A _5196_/B _5196_/C vssd1 vssd1 vccd1 vccd1 _5242_/B sky130_fd_sc_hd__a21oi_1
X_6488__70 vssd1 vssd1 vccd1 vccd1 _6488__70/HI _6596_/A sky130_fd_sc_hd__conb_1
X_5172_ _5172_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5208_/B sky130_fd_sc_hd__xnor2_2
X_4123_ _4122_/B _4122_/C _4122_/D _4122_/A vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__o22a_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4054_ _5159_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4956_ _4956_/A _4956_/B vssd1 vssd1 vccd1 vccd1 _4957_/A sky130_fd_sc_hd__nand2_1
X_3907_ _5424_/A vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__buf_2
X_4887_ _4895_/C vssd1 vssd1 vccd1 vccd1 _4956_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6626_ _6626_/A _3324_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_3838_ _3854_/A _3854_/B vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__nand2_1
X_6557_ _6557_/A _3243_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3769_ _3871_/A _3871_/B _3604_/A vssd1 vssd1 vccd1 vccd1 _3813_/B sky130_fd_sc_hd__a21o_2
X_5508_ _5508_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__xnor2_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5439_ _5362_/A _5350_/B _5467_/A vssd1 vssd1 vccd1 vccd1 _5439_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4810_ _4810_/A _4810_/B vssd1 vssd1 vccd1 vccd1 _4811_/B sky130_fd_sc_hd__xnor2_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5790_ _5790_/A _5790_/B vssd1 vssd1 vccd1 vccd1 _5790_/Y sky130_fd_sc_hd__xnor2_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4939_/A _4939_/B vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__xnor2_1
X_4672_ _6060_/A _3566_/A _4648_/B _4642_/D vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__o31a_1
X_3623_ _3624_/A _3651_/A vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__and2_1
X_6411_ _6426_/CLK _6411_/D vssd1 vssd1 vccd1 vccd1 _6411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3554_ _3554_/A _3554_/B vssd1 vssd1 vccd1 vccd1 _3585_/B sky130_fd_sc_hd__nand2_1
X_6342_ _6345_/CLK _6342_/D vssd1 vssd1 vccd1 vccd1 _6342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3485_ _3485_/A _3485_/B vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__xnor2_1
X_6273_ _6273_/A _6294_/B vssd1 vssd1 vccd1 vccd1 _6410_/D sky130_fd_sc_hd__nor2_1
X_5224_ _5221_/X _5222_/X _5225_/A _5223_/X vssd1 vssd1 vccd1 vccd1 _5225_/B sky130_fd_sc_hd__a211oi_2
XFILLER_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5155_ _5155_/A _5155_/B vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4106_ _4298_/B vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__clkbuf_2
X_5086_ _5592_/A _5592_/B vssd1 vssd1 vccd1 vccd1 _5090_/C sky130_fd_sc_hd__nor2_1
X_4037_ _4037_/A vssd1 vssd1 vccd1 vccd1 _4037_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5988_ _6014_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _5988_/Y sky130_fd_sc_hd__nand2_1
X_4939_ _4939_/A _4939_/B vssd1 vssd1 vccd1 vccd1 _4939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6609_ _6609_/A _3314_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _3272_/A vssd1 vssd1 vccd1 vccd1 _3270_/Y sky130_fd_sc_hd__inv_2
X_6458__40 vssd1 vssd1 vccd1 vccd1 _6458__40/HI _6563_/A sky130_fd_sc_hd__conb_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5911_ _6100_/A vssd1 vssd1 vccd1 vccd1 _5911_/X sky130_fd_sc_hd__clkbuf_4
X_5842_ _5842_/A vssd1 vssd1 vccd1 vccd1 _5945_/A sky130_fd_sc_hd__buf_2
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5773_ _5783_/A _5783_/B vssd1 vssd1 vccd1 vccd1 _5784_/B sky130_fd_sc_hd__nor2_1
X_4724_ _4724_/A _4724_/B vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__or2_1
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4655_ _4655_/A _4655_/B vssd1 vssd1 vccd1 vccd1 _4655_/Y sky130_fd_sc_hd__nor2_1
X_3606_ _6330_/Q vssd1 vssd1 vccd1 vccd1 _5997_/A sky130_fd_sc_hd__inv_2
X_4586_ _5067_/A _4586_/B vssd1 vssd1 vccd1 vccd1 _4586_/X sky130_fd_sc_hd__or2_1
X_6325_ _6426_/CLK _6325_/D vssd1 vssd1 vccd1 vccd1 _6325_/Q sky130_fd_sc_hd__dfxtp_1
X_3537_ _4642_/D vssd1 vssd1 vccd1 vccd1 _4694_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3468_ _3469_/B _3469_/C _3469_/A vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__a21oi_1
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6256_ _6404_/Q _6403_/Q _6256_/C vssd1 vssd1 vccd1 vccd1 _6262_/C sky130_fd_sc_hd__and3_1
X_5207_ _5207_/A _5253_/A vssd1 vssd1 vccd1 vccd1 _5210_/A sky130_fd_sc_hd__or2_2
X_3399_ _4765_/D vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6187_ _6187_/A vssd1 vssd1 vccd1 vccd1 _6377_/D sky130_fd_sc_hd__clkbuf_1
X_5138_ _5711_/A _5029_/B _5125_/B _5137_/Y vssd1 vssd1 vccd1 vccd1 _5144_/B sky130_fd_sc_hd__a31oi_2
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5069_ _5137_/B _5070_/B vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__or2_1
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4573_/A _4573_/B _4440_/C vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__or3_1
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4371_ _5471_/C _4393_/B vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__and2_1
X_6110_ _6347_/Q _6115_/B vssd1 vssd1 vccd1 vccd1 _6111_/A sky130_fd_sc_hd__and2_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3322_ _3334_/A vssd1 vssd1 vccd1 vccd1 _3327_/A sky130_fd_sc_hd__buf_12
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3253_ _3253_/A vssd1 vssd1 vccd1 vccd1 _3253_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6041_/A vssd1 vssd1 vccd1 vccd1 _6099_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5825_ _5825_/A vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5756_ _5756_/A _5978_/A _5756_/C _5756_/D vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__or4_4
X_4707_ _4701_/A _4701_/B _4706_/X vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__o21ba_1
X_5687_ _5688_/A _5688_/B vssd1 vssd1 vccd1 vccd1 _5691_/B sky130_fd_sc_hd__xor2_1
X_4638_ _5823_/B vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4569_ _4569_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6308_ _6423_/Q _6309_/C _6307_/Y vssd1 vssd1 vccd1 vccd1 _6423_/D sky130_fd_sc_hd__o21a_1
X_6239_ _6397_/Q _6243_/B vssd1 vssd1 vccd1 vccd1 _6240_/A sky130_fd_sc_hd__and2_1
XFILLER_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6428__10 vssd1 vssd1 vccd1 vccd1 _6428__10/HI _6533_/A sky130_fd_sc_hd__conb_1
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3940_ _4317_/B vssd1 vssd1 vccd1 vccd1 _4302_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3871_ _3871_/A _3871_/B vssd1 vssd1 vccd1 vccd1 _4068_/B sky130_fd_sc_hd__xor2_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6590_ _6590_/A _3282_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
X_5610_ _5091_/A _5054_/B _5054_/A vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__o21ba_1
X_5541_ _5543_/A _5543_/B vssd1 vssd1 vccd1 vccd1 _5568_/B sky130_fd_sc_hd__or2_1
XFILLER_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5472_ _5473_/A _5500_/A vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__nand2_1
X_4423_ _6316_/Q vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4354_ _4354_/A _4354_/B vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__xor2_1
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3305_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4285_ _4305_/A _4284_/Y _4284_/A vssd1 vssd1 vccd1 vccd1 _4290_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6024_ _6024_/A vssd1 vssd1 vccd1 vccd1 _6334_/D sky130_fd_sc_hd__clkbuf_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3248_/A vssd1 vssd1 vccd1 vccd1 _3241_/A sky130_fd_sc_hd__buf_12
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5808_ _5842_/A _5746_/X _5806_/X _5807_/X vssd1 vssd1 vccd1 vccd1 _5808_/Y sky130_fd_sc_hd__a22oi_2
X_5739_ _5766_/B _5775_/A _5787_/A _5758_/A _5766_/A vssd1 vssd1 vccd1 vccd1 _5796_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6512__94 vssd1 vssd1 vccd1 vccd1 _6512__94/HI _6620_/A sky130_fd_sc_hd__conb_1
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _4069_/A _4069_/B _5248_/B _4152_/B vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4972_ _4948_/A _4967_/B _4948_/C _4793_/X vssd1 vssd1 vccd1 vccd1 _4973_/B sky130_fd_sc_hd__a31o_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _3921_/A _3921_/B _3922_/X vssd1 vssd1 vccd1 vccd1 _4476_/B sky130_fd_sc_hd__a21bo_1
XFILLER_32_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3854_ _3854_/A _3854_/B vssd1 vssd1 vccd1 vccd1 _3855_/B sky130_fd_sc_hd__or2_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3785_ _3960_/A vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__buf_2
X_6573_ _6573_/A _3262_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5524_ _5524_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _5524_/Y sky130_fd_sc_hd__nor2_1
X_5455_ _5545_/A _5455_/B _5455_/C vssd1 vssd1 vccd1 vccd1 _5476_/A sky130_fd_sc_hd__and3_1
X_4406_ _5518_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4424_/C sky130_fd_sc_hd__and2_1
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5386_ _5386_/A _5492_/B _5492_/C vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__and3_1
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4337_ _4307_/A _4436_/B _4272_/B vssd1 vssd1 vccd1 vccd1 _4338_/B sky130_fd_sc_hd__a21oi_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _4268_/A _4268_/B vssd1 vssd1 vccd1 vccd1 _4279_/B sky130_fd_sc_hd__or2_1
X_6007_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6007_/X sky130_fd_sc_hd__buf_4
X_3219_ _3222_/A vssd1 vssd1 vccd1 vccd1 _3219_/Y sky130_fd_sc_hd__inv_2
X_4199_ _4199_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4246_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3647_/A _3646_/C _3570_/C vssd1 vssd1 vccd1 vccd1 _3570_/X sky130_fd_sc_hd__and3_1
XFILLER_115_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5240_ _5281_/A _5240_/B _5240_/C vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__and3_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5171_ _5178_/A _5212_/A _5170_/X vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__o21a_1
X_4122_ _4122_/A _4122_/B _4122_/C _4122_/D vssd1 vssd1 vccd1 vccd1 _4122_/Y sky130_fd_sc_hd__nor4_2
X_4053_ _4037_/A _4025_/B _4025_/C vssd1 vssd1 vccd1 vccd1 _4075_/B sky130_fd_sc_hd__a21o_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4955_ _5275_/A _4955_/B vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__xor2_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3906_ _5486_/A vssd1 vssd1 vccd1 vccd1 _5424_/A sky130_fd_sc_hd__clkbuf_2
X_4886_ _4886_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _4886_/Y sky130_fd_sc_hd__nand2_1
X_6625_ _6625_/A _3323_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_3837_ _3837_/A _3857_/A vssd1 vssd1 vccd1 vccd1 _3854_/B sky130_fd_sc_hd__or2_1
X_3768_ _3894_/A _3894_/B _3767_/Y vssd1 vssd1 vccd1 vccd1 _3871_/B sky130_fd_sc_hd__a21o_2
X_6556_ _6556_/A _3241_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_5507_ _5509_/A _5509_/B _5506_/X vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__a21bo_2
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3699_ _3699_/A _4895_/B _3699_/C _3699_/D vssd1 vssd1 vccd1 vccd1 _3726_/A sky130_fd_sc_hd__and4_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5438_ _5467_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5438_/X sky130_fd_sc_hd__and2b_1
X_5369_ _5369_/A _5369_/B vssd1 vssd1 vccd1 vccd1 _5487_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4740_/A _4740_/B vssd1 vssd1 vccd1 vccd1 _4939_/B sky130_fd_sc_hd__nor2_1
X_4671_ _6340_/Q vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__clkbuf_2
X_3622_ _3685_/A _3650_/B _4800_/C vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__a21o_1
X_6410_ _6426_/CLK _6410_/D vssd1 vssd1 vccd1 vccd1 _6410_/Q sky130_fd_sc_hd__dfxtp_1
X_6341_ _6345_/CLK _6341_/D vssd1 vssd1 vccd1 vccd1 _6341_/Q sky130_fd_sc_hd__dfxtp_1
X_3553_ _3553_/A _3553_/B _3553_/C vssd1 vssd1 vccd1 vccd1 _3554_/B sky130_fd_sc_hd__nand3_1
X_3484_ _3484_/A _3484_/B vssd1 vssd1 vccd1 vccd1 _3516_/A sky130_fd_sc_hd__xor2_1
X_6272_ _6409_/Q _6269_/B _6271_/Y vssd1 vssd1 vccd1 vccd1 _6409_/D sky130_fd_sc_hd__o21a_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5223_ _5219_/X _5218_/Y _5217_/X _5209_/Y vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__o211a_1
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _5154_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5155_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4105_ _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4298_/B sky130_fd_sc_hd__and2_1
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5085_ _5085_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5592_/B sky130_fd_sc_hd__xnor2_1
X_4036_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5712_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5987_ _5987_/A _5987_/B vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__xnor2_1
X_4938_ _4974_/A _4974_/B _4977_/B vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__or3_1
X_4869_ _4859_/A _4858_/B _4858_/C vssd1 vssd1 vccd1 vccd1 _4878_/B sky130_fd_sc_hd__a21o_1
X_6608_ _6608_/A _3339_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539_ _6539_/A _3220_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6473__55 vssd1 vssd1 vccd1 vccd1 _6473__55/HI _6581_/A sky130_fd_sc_hd__conb_1
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _6025_/B vssd1 vssd1 vccd1 vccd1 _6100_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5841_ _6413_/Q _5827_/X _5840_/Y _6414_/Q vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__o22a_1
X_5772_ _5765_/X _5746_/X _5770_/X _5807_/A vssd1 vssd1 vccd1 vccd1 _5783_/B sky130_fd_sc_hd__a22o_1
X_4723_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__or2_1
X_4654_ _4655_/A _4655_/B vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__xor2_1
X_3605_ _3605_/A _3605_/B vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__xnor2_4
X_4585_ _4571_/X _4583_/X _4584_/X vssd1 vssd1 vccd1 vccd1 _4588_/B sky130_fd_sc_hd__o21ai_1
X_6324_ _6388_/CLK _6324_/D vssd1 vssd1 vccd1 vccd1 _6324_/Q sky130_fd_sc_hd__dfxtp_1
X_3536_ _6328_/Q _4642_/D _3538_/C _6326_/Q vssd1 vssd1 vccd1 vccd1 _3547_/A sky130_fd_sc_hd__a22o_2
X_6255_ _6403_/Q _6256_/C _6404_/Q vssd1 vssd1 vccd1 vccd1 _6257_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3467_ _3467_/A _3467_/B vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5206_ _5252_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _5253_/A sky130_fd_sc_hd__and2_1
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3398_ _3653_/A vssd1 vssd1 vccd1 vccd1 _4765_/D sky130_fd_sc_hd__buf_2
X_6186_ _6376_/Q _6194_/B vssd1 vssd1 vccd1 vccd1 _6187_/A sky130_fd_sc_hd__and2_1
X_5137_ _5137_/A _5137_/B vssd1 vssd1 vccd1 vccd1 _5137_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5068_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5070_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4019_ _5281_/A _4068_/B vssd1 vssd1 vccd1 vccd1 _4021_/C sky130_fd_sc_hd__and2_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4370_ _4370_/A _4370_/B vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__xor2_1
X_3321_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3321_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3252_ _3253_/A vssd1 vssd1 vccd1 vccd1 _3252_/Y sky130_fd_sc_hd__inv_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6040_/B vssd1 vssd1 vccd1 vccd1 _6040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5824_ _5807_/X _5821_/X _5825_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5824_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5755_ _5979_/A vssd1 vssd1 vccd1 vccd1 _5978_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4706_ _4702_/B _4706_/B vssd1 vssd1 vccd1 vccd1 _4706_/X sky130_fd_sc_hd__and2b_1
X_5686_ _5686_/A _5686_/B vssd1 vssd1 vccd1 vccd1 _5688_/B sky130_fd_sc_hd__nand2_1
X_4637_ _5871_/A _6103_/A _5817_/A vssd1 vssd1 vccd1 vccd1 _5823_/B sky130_fd_sc_hd__nor3_2
X_4568_ _4569_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4571_/B sky130_fd_sc_hd__xor2_1
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ _3519_/A _3519_/B vssd1 vssd1 vccd1 vccd1 _3520_/B sky130_fd_sc_hd__nand2_1
X_6307_ _6310_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6307_/Y sky130_fd_sc_hd__nor2_1
X_4499_ _4499_/A vssd1 vssd1 vccd1 vccd1 _4499_/Y sky130_fd_sc_hd__inv_2
X_6238_ _6238_/A vssd1 vssd1 vccd1 vccd1 _6397_/D sky130_fd_sc_hd__clkbuf_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6370_/Q _6183_/B vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__and2_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6443__25 vssd1 vssd1 vccd1 vccd1 _6443__25/HI _6548_/A sky130_fd_sc_hd__conb_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _3870_/A _3870_/B vssd1 vssd1 vccd1 vccd1 _3879_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5540_ _5544_/A _5544_/B _5537_/A vssd1 vssd1 vccd1 vccd1 _5543_/B sky130_fd_sc_hd__o21ba_1
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5471_ _5471_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5500_/A sky130_fd_sc_hd__and3_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4422_ _4422_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4448_/A sky130_fd_sc_hd__xnor2_1
X_4353_ _4459_/B _4353_/B vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__xnor2_4
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4284_ _4284_/A _4284_/B vssd1 vssd1 vccd1 vccd1 _4284_/Y sky130_fd_sc_hd__nor2_1
X_3304_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__buf_8
X_3235_ _3235_/A vssd1 vssd1 vccd1 vccd1 _3235_/Y sky130_fd_sc_hd__inv_2
X_6023_ _6392_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6024_/A sky130_fd_sc_hd__and2_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3999_ _3980_/Y _3996_/X _3997_/X _3998_/Y vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__a211oi_2
X_5807_ _5807_/A vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__buf_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5738_ _5738_/A vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__inv_2
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5669_/A _5709_/A vssd1 vssd1 vccd1 vccd1 _5726_/A sky130_fd_sc_hd__xnor2_1
XFILLER_116_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4971_ _4971_/A _4971_/B vssd1 vssd1 vccd1 vccd1 _4973_/A sky130_fd_sc_hd__nand2_1
X_3922_ _3953_/A _3953_/B vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__or2b_1
X_3853_ _3887_/A _3853_/B vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__xor2_4
XFILLER_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3784_ _5282_/A vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__clkbuf_2
X_6572_ _6572_/A _3260_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5523_ _5530_/A _5523_/B vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__and2_1
XFILLER_117_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5454_ _5454_/A _5454_/B vssd1 vssd1 vccd1 vccd1 _5484_/A sky130_fd_sc_hd__xnor2_4
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5385_ _5385_/A _5385_/B vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__xnor2_4
X_4405_ _5967_/A _5486_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _5545_/C sky130_fd_sc_hd__and3_1
X_4336_ _4336_/A vssd1 vssd1 vccd1 vccd1 _4436_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _4307_/A _4406_/B _4235_/C vssd1 vssd1 vccd1 vccd1 _4268_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4198_ _4208_/A _4208_/B vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__and2_1
X_3218_ _3222_/A vssd1 vssd1 vccd1 vccd1 _3218_/Y sky130_fd_sc_hd__inv_2
X_6006_ _5992_/X _6004_/X _6005_/Y _6014_/A vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__o211a_1
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5170_ _5096_/A _5101_/B _5096_/B _5095_/A vssd1 vssd1 vccd1 vccd1 _5170_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4121_ _4121_/A _4121_/B _4121_/C _4121_/D vssd1 vssd1 vccd1 vccd1 _4121_/Y sky130_fd_sc_hd__nand4_4
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4052_ _4050_/A _4049_/C _4049_/B vssd1 vssd1 vccd1 vccd1 _4472_/B sky130_fd_sc_hd__a21o_1
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _4953_/A _4953_/B _4953_/C vssd1 vssd1 vccd1 vccd1 _5231_/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3905_ _6318_/Q vssd1 vssd1 vccd1 vccd1 _5486_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _4885_/A _4885_/B vssd1 vssd1 vccd1 vccd1 _4907_/A sky130_fd_sc_hd__xnor2_1
X_3836_ _3856_/A _3856_/B vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__and2_1
X_6624_ _6624_/A _3321_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
X_3767_ _3767_/A _3767_/B vssd1 vssd1 vccd1 vccd1 _3767_/Y sky130_fd_sc_hd__nor2_1
X_6555_ _6555_/A _3240_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
X_5506_ _5506_/A _5505_/A vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__or2b_1
X_3698_ _3692_/A _3691_/C _3691_/B vssd1 vssd1 vccd1 vccd1 _3707_/B sky130_fd_sc_hd__a21o_1
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5437_ _5390_/B _5475_/A _5426_/X vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__a21bo_1
X_5368_ _5368_/A _5368_/B vssd1 vssd1 vccd1 vccd1 _5369_/B sky130_fd_sc_hd__or2_1
X_6479__61 vssd1 vssd1 vccd1 vccd1 _6479__61/HI _6587_/A sky130_fd_sc_hd__conb_1
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4327_/A _4327_/B vssd1 vssd1 vccd1 vccd1 _4349_/B sky130_fd_sc_hd__xor2_1
XFILLER_87_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5299_ _5335_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5305_/B sky130_fd_sc_hd__and2_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6526__108 vssd1 vssd1 vccd1 vccd1 _6526__108/HI _6634_/A sky130_fd_sc_hd__conb_1
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4765_/D _4802_/B vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__nand2_1
X_3621_ _6332_/Q _4805_/B vssd1 vssd1 vccd1 vccd1 _4800_/C sky130_fd_sc_hd__and2_1
X_3552_ _3553_/B _3553_/C _3553_/A vssd1 vssd1 vccd1 vccd1 _3554_/A sky130_fd_sc_hd__a21o_1
X_6340_ _6345_/CLK _6340_/D vssd1 vssd1 vccd1 vccd1 _6340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3483_ _3483_/A _3518_/A _3482_/X vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__or3b_1
X_6271_ _6409_/Q _6269_/B _6007_/X vssd1 vssd1 vccd1 vccd1 _6271_/Y sky130_fd_sc_hd__a21oi_1
X_5222_ _5222_/A _5216_/B vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__or2b_1
XFILLER_69_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5153_ _5153_/A _5153_/B vssd1 vssd1 vccd1 vccd1 _5188_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ _4104_/A _4213_/D _4135_/A vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__and3_1
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5084_ _5085_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5090_/B sky130_fd_sc_hd__and2_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _5257_/A vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__buf_2
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _5967_/A _5980_/B _5978_/X vssd1 vssd1 vccd1 vccd1 _5987_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _4937_/A _4937_/B vssd1 vssd1 vccd1 vccd1 _4977_/B sky130_fd_sc_hd__xnor2_4
X_4868_ _4866_/A _4864_/Y _4862_/X _4863_/X vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__o211a_1
X_6607_ _6607_/A _3302_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
X_3819_ _3808_/A _3875_/A _3817_/Y _3870_/A vssd1 vssd1 vccd1 vccd1 _3835_/B sky130_fd_sc_hd__o22a_1
X_4799_ _4805_/A _4805_/C _4830_/D _4805_/B vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__or4b_1
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6538_ _6538_/A _3219_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5840_ _5936_/A _5825_/X _5839_/X _5807_/X vssd1 vssd1 vccd1 vccd1 _5840_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ _5771_/A vssd1 vssd1 vccd1 vccd1 _5807_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4722_ _4722_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__or2_1
X_4653_ _4886_/A _4749_/B vssd1 vssd1 vccd1 vccd1 _4655_/B sky130_fd_sc_hd__nand2_1
X_3604_ _3604_/A _3604_/B vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__nor2_2
X_4584_ _5711_/A _4580_/X _4583_/B _4583_/A vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__a211o_1
X_3535_ _3535_/A _3576_/A vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__xnor2_2
X_6323_ _6361_/CLK _6323_/D vssd1 vssd1 vccd1 vccd1 _6323_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3466_ _3466_/A _3466_/B _3466_/C vssd1 vssd1 vccd1 vccd1 _3467_/B sky130_fd_sc_hd__nand3_1
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6254_ _6403_/Q _6256_/C _6253_/Y vssd1 vssd1 vccd1 vccd1 _6403_/D sky130_fd_sc_hd__o21a_1
X_6449__31 vssd1 vssd1 vccd1 vccd1 _6449__31/HI _6554_/A sky130_fd_sc_hd__conb_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5205_ _5205_/A _5205_/B vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__xnor2_1
X_3397_ _3592_/D vssd1 vssd1 vccd1 vccd1 _3406_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6185_ _6234_/A vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5136_ _5136_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5144_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5067_ _5067_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5137_/B sky130_fd_sc_hd__nand2_1
X_4018_ _4989_/A _4302_/B _4055_/B _4016_/Y vssd1 vssd1 vccd1 vccd1 _4024_/B sky130_fd_sc_hd__a31o_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5969_ _6324_/Q _6335_/Q vssd1 vssd1 vccd1 vccd1 _5969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3320_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3320_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3253_/A vssd1 vssd1 vccd1 vccd1 _3251_/Y sky130_fd_sc_hd__inv_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5823_ _5868_/A _5823_/B _5823_/C vssd1 vssd1 vccd1 vccd1 _5825_/A sky130_fd_sc_hd__or3_1
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5754_ _6408_/Q _5753_/X _5744_/X _6409_/Q vssd1 vssd1 vccd1 vccd1 _5754_/X sky130_fd_sc_hd__o22a_1
X_4705_ _4791_/A _4791_/B _4704_/X vssd1 vssd1 vccd1 vccd1 _4919_/A sky130_fd_sc_hd__a21bo_1
X_5685_ _5693_/A _5699_/A _5564_/B vssd1 vssd1 vccd1 vccd1 _5686_/B sky130_fd_sc_hd__a21o_1
X_4636_ _4636_/A vssd1 vssd1 vccd1 vccd1 _6103_/A sky130_fd_sc_hd__buf_2
X_4567_ _4567_/A _4567_/B vssd1 vssd1 vccd1 vccd1 _4569_/B sky130_fd_sc_hd__nand2_1
X_6306_ _6423_/Q _6309_/C vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__and2_1
X_3518_ _3518_/A _3518_/B _3561_/A vssd1 vssd1 vccd1 vccd1 _3804_/B sky130_fd_sc_hd__nand3_1
X_4498_ _4498_/A vssd1 vssd1 vccd1 vccd1 _4498_/Y sky130_fd_sc_hd__inv_2
X_3449_ _3449_/A _3449_/B vssd1 vssd1 vccd1 vccd1 _3463_/A sky130_fd_sc_hd__nor2_1
X_6237_ _6396_/Q _6243_/B vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__and2_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6168_/A vssd1 vssd1 vccd1 vccd1 _6370_/D sky130_fd_sc_hd__clkbuf_1
X_5119_ _5119_/A _5119_/B vssd1 vssd1 vccd1 vccd1 _5132_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6099_ _6099_/A _6099_/B vssd1 vssd1 vccd1 vccd1 _6099_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6361_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5470_ _5470_/A _5470_/B vssd1 vssd1 vccd1 vccd1 _5473_/A sky130_fd_sc_hd__xnor2_1
XFILLER_117_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4421_ _4421_/A _4453_/A vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__xor2_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4352_ _4321_/B _4328_/X _4350_/B _4351_/Y vssd1 vssd1 vccd1 vccd1 _4353_/B sky130_fd_sc_hd__o31a_2
X_4283_ _4304_/A _4304_/B vssd1 vssd1 vccd1 vccd1 _4284_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3303_ _3303_/A vssd1 vssd1 vccd1 vccd1 _3303_/Y sky130_fd_sc_hd__inv_2
X_3234_ _3235_/A vssd1 vssd1 vccd1 vccd1 _3234_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6022_/A vssd1 vssd1 vccd1 vccd1 _6333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3998_ _3997_/A _3997_/C _3997_/B vssd1 vssd1 vccd1 vccd1 _3998_/Y sky130_fd_sc_hd__a21oi_2
X_5806_ _4639_/A _5804_/X _5805_/X _5868_/B vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5737_ _5774_/A _5774_/B _5774_/C vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__a21oi_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5668_ _5727_/A _5727_/B vssd1 vssd1 vccd1 vccd1 _5668_/X sky130_fd_sc_hd__or2_1
X_4619_ _5750_/A _5805_/A _5805_/B _4618_/Y vssd1 vssd1 vccd1 vccd1 _4619_/X sky130_fd_sc_hd__a31o_1
X_5599_ _5613_/A _5613_/B _5091_/A vssd1 vssd1 vccd1 vccd1 _5600_/B sky130_fd_sc_hd__a21o_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6503__85 vssd1 vssd1 vccd1 vccd1 _6503__85/HI _6611_/A sky130_fd_sc_hd__conb_1
XFILLER_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4970_ _4970_/A _4970_/B vssd1 vssd1 vccd1 vccd1 _4971_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3921_ _3921_/A _3921_/B vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__xor2_1
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3852_ _3887_/B _3852_/B vssd1 vssd1 vccd1 vccd1 _3853_/B sky130_fd_sc_hd__xnor2_2
X_6571_ _6571_/A _3259_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
X_3783_ _5237_/A vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__clkbuf_2
X_5522_ _4373_/A _5236_/A _5511_/Y _5514_/X vssd1 vssd1 vccd1 vccd1 _5523_/B sky130_fd_sc_hd__a211o_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5453_ _5453_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _5655_/A sky130_fd_sc_hd__xnor2_2
X_5384_ _5580_/B _5384_/B vssd1 vssd1 vccd1 vccd1 _5636_/A sky130_fd_sc_hd__xnor2_4
X_4404_ _4404_/A vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__buf_2
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4335_ _4335_/A _4335_/B vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4266_ _4266_/A _4266_/B vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4197_ _4199_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__and2_1
X_3217_ _3342_/A vssd1 vssd1 vccd1 vccd1 _3222_/A sky130_fd_sc_hd__clkbuf_16
X_6005_ _4629_/B _5998_/X _5992_/X vssd1 vssd1 vccd1 vccd1 _6005_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4120_ _4113_/A _4113_/B _4113_/C vssd1 vssd1 vccd1 vccd1 _4121_/D sky130_fd_sc_hd__o21ai_2
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4051_ _4474_/A _4474_/B _4474_/C vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4953_ _4953_/A _4953_/B _4953_/C vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__and3_1
X_3904_ _5122_/A _3903_/B _3903_/C vssd1 vssd1 vccd1 vccd1 _3915_/B sky130_fd_sc_hd__a21oi_1
X_6623_ _6623_/A _3320_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4884_ _4882_/A _4882_/C _4882_/B vssd1 vssd1 vccd1 vccd1 _4909_/B sky130_fd_sc_hd__a21o_1
X_3835_ _3835_/A _3835_/B vssd1 vssd1 vccd1 vccd1 _3856_/B sky130_fd_sc_hd__xnor2_1
X_6554_ _6554_/A _3239_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
X_3766_ _3938_/A _3938_/B _3765_/X vssd1 vssd1 vccd1 vccd1 _3894_/B sky130_fd_sc_hd__a21o_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5505_ _5505_/A _5506_/A vssd1 vssd1 vccd1 vccd1 _5509_/B sky130_fd_sc_hd__xnor2_1
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3697_ _3697_/A _3697_/B vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__xnor2_4
X_5436_ _5436_/A _5436_/B vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _5367_/A _5546_/B vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__nand2_1
X_4318_ _4318_/A _4318_/B vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__xor2_2
X_5298_ _5289_/A _5289_/B _5297_/X vssd1 vssd1 vccd1 vccd1 _5300_/A sky130_fd_sc_hd__o21ba_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4201_/B _4209_/X _4247_/B _4248_/X vssd1 vssd1 vccd1 vccd1 _4250_/B sky130_fd_sc_hd__a31oi_4
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6494__76 vssd1 vssd1 vccd1 vccd1 _6494__76/HI _6602_/A sky130_fd_sc_hd__conb_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _3671_/B vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3551_ _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3553_/A sky130_fd_sc_hd__nand2_1
X_3482_ _3482_/A _3482_/B vssd1 vssd1 vccd1 vccd1 _3482_/X sky130_fd_sc_hd__and2_1
X_6270_ _6408_/Q _6266_/B _6269_/Y vssd1 vssd1 vccd1 vccd1 _6408_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5221_ _5221_/A _5215_/A vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__or2b_1
X_5152_ _5152_/A _5152_/B vssd1 vssd1 vccd1 vccd1 _5153_/B sky130_fd_sc_hd__or2_1
XFILLER_69_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4103_ _5371_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__and3_1
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5083_ _5083_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _5085_/B sky130_fd_sc_hd__xor2_1
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4034_ _5335_/A vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _5985_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__xnor2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _4941_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__and2b_1
X_4867_ _4913_/B _4867_/B vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__xnor2_4
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _3818_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__nand2_1
X_6606_ _6606_/A _3301_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_4798_ _4798_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__or2_1
X_6537_ _6537_/A _3218_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_3749_ _4886_/B vssd1 vssd1 vccd1 vccd1 _4577_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5419_ _5418_/B _5419_/B vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__and2b_1
X_6399_ _6401_/CLK _6399_/D vssd1 vssd1 vccd1 vccd1 _6399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5770_ _4639_/A _5767_/X _5769_/Y _5868_/B vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__a22o_1
X_4721_ _4919_/A _4919_/B vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__and2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4652_ _6342_/Q _3473_/B _4751_/C vssd1 vssd1 vccd1 vccd1 _4749_/B sky130_fd_sc_hd__mux2_2
X_3603_ _3603_/A _3603_/B vssd1 vssd1 vccd1 vccd1 _3604_/B sky130_fd_sc_hd__and2_1
X_4583_ _4583_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4583_/X sky130_fd_sc_hd__and2_1
XFILLER_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3534_ _4677_/A _4888_/A _3716_/C _3534_/D vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__and4_2
X_6322_ _6361_/CLK _6322_/D vssd1 vssd1 vccd1 vccd1 _6322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3465_ _3485_/A _3485_/B vssd1 vssd1 vccd1 vccd1 _3469_/C sky130_fd_sc_hd__or2_1
X_6253_ _6403_/Q _6256_/C _6007_/X vssd1 vssd1 vccd1 vccd1 _6253_/Y sky130_fd_sc_hd__a21oi_1
X_5204_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5205_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3396_ _3406_/C _6010_/A _3407_/A vssd1 vssd1 vccd1 vccd1 _3441_/A sky130_fd_sc_hd__mux2_1
X_6184_ _6184_/A vssd1 vssd1 vccd1 vccd1 _6376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5135_ _5145_/A _5135_/B vssd1 vssd1 vccd1 vccd1 _5140_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6464__46 vssd1 vssd1 vccd1 vccd1 _6464__46/HI _6569_/A sky130_fd_sc_hd__conb_1
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ _5072_/A _5072_/B vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__xnor2_1
X_4017_ _3966_/B _4014_/Y _4016_/Y vssd1 vssd1 vccd1 vccd1 _4055_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5968_ _6324_/Q _6335_/Q vssd1 vssd1 vccd1 vccd1 _5968_/X sky130_fd_sc_hd__and2_1
X_4919_ _4919_/A _4919_/B vssd1 vssd1 vccd1 vccd1 _4970_/B sky130_fd_sc_hd__xor2_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5899_ _6425_/Q _5896_/B _6310_/A vssd1 vssd1 vccd1 vccd1 _5899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3253_/A vssd1 vssd1 vccd1 vccd1 _3250_/Y sky130_fd_sc_hd__inv_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5822_ _6106_/A _6103_/A _5848_/A vssd1 vssd1 vccd1 vccd1 _5823_/C sky130_fd_sc_hd__and3b_1
X_5753_ _5851_/A _5746_/X _5752_/X _4634_/X vssd1 vssd1 vccd1 vccd1 _5753_/X sky130_fd_sc_hd__o2bb2a_1
X_4704_ _4704_/A _4703_/B vssd1 vssd1 vccd1 vccd1 _4704_/X sky130_fd_sc_hd__or2b_1
X_5684_ _5684_/A _5684_/B vssd1 vssd1 vccd1 vccd1 _5723_/A sky130_fd_sc_hd__xnor2_1
X_6509__91 vssd1 vssd1 vccd1 vccd1 _6509__91/HI _6617_/A sky130_fd_sc_hd__conb_1
X_4635_ _3354_/X _5745_/B _4619_/X _5868_/B _4634_/X vssd1 vssd1 vccd1 vccd1 _4635_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _4575_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4567_/B sky130_fd_sc_hd__nand2_1
X_3517_ _3560_/A _3560_/B vssd1 vssd1 vccd1 vccd1 _3561_/A sky130_fd_sc_hd__or2_1
X_6305_ _6422_/Q _6301_/B _6304_/Y vssd1 vssd1 vccd1 vccd1 _6422_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4497_ _4497_/A _4497_/B vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__xor2_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3448_ _4886_/A _3395_/B _3430_/C vssd1 vssd1 vccd1 vccd1 _3449_/B sky130_fd_sc_hd__a21oi_1
X_6236_ _6236_/A vssd1 vssd1 vccd1 vccd1 _6396_/D sky130_fd_sc_hd__clkbuf_1
X_3379_ _3395_/A vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__clkbuf_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6369_/Q _6183_/B vssd1 vssd1 vccd1 vccd1 _6168_/A sky130_fd_sc_hd__and2_1
X_5118_ _5118_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6098_ _6097_/A _6103_/C _6097_/C vssd1 vssd1 vccd1 vccd1 _6099_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5049_ _5602_/A _5049_/B vssd1 vssd1 vccd1 vccd1 _5050_/B sky130_fd_sc_hd__and2_1
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4420_ _4451_/A _4451_/B _4419_/A vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__a21oi_2
XFILLER_113_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4351_ _4354_/A _4354_/B vssd1 vssd1 vccd1 vccd1 _4351_/Y sky130_fd_sc_hd__nand2_1
X_4282_ _4304_/A _4304_/B vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__and2_1
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3302_ _3303_/A vssd1 vssd1 vccd1 vccd1 _3302_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3233_ _3235_/A vssd1 vssd1 vccd1 vccd1 _3233_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6019_/X _6021_/B vssd1 vssd1 vccd1 vccd1 _6022_/A sky130_fd_sc_hd__and2b_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6434__16 vssd1 vssd1 vccd1 vccd1 _6434__16/HI _6539_/A sky130_fd_sc_hd__conb_1
XFILLER_94_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3997_ _3997_/A _3997_/B _3997_/C vssd1 vssd1 vccd1 vccd1 _3997_/X sky130_fd_sc_hd__and3_1
X_5805_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5805_/X sky130_fd_sc_hd__xor2_2
X_5736_ _5736_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _5774_/C sky130_fd_sc_hd__xnor2_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _5672_/A _5665_/X _5671_/A vssd1 vssd1 vccd1 vccd1 _5727_/B sky130_fd_sc_hd__a21oi_1
X_4618_ _4618_/A vssd1 vssd1 vccd1 vccd1 _4618_/Y sky130_fd_sc_hd__inv_2
X_5598_ _5654_/A _5654_/B _5639_/A _5597_/Y vssd1 vssd1 vccd1 vccd1 _5613_/B sky130_fd_sc_hd__a31o_2
X_4549_ _4549_/A _4549_/B vssd1 vssd1 vccd1 vccd1 _4549_/X sky130_fd_sc_hd__or2_1
XFILLER_8_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6219_ _6219_/A vssd1 vssd1 vccd1 vccd1 _6390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3920_ _3915_/A _3920_/B vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__and2b_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3851_ _3844_/A _3849_/Y _4499_/A vssd1 vssd1 vccd1 vccd1 _3852_/B sky130_fd_sc_hd__a21o_1
X_6570_ _6570_/A _3258_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_3782_ _5316_/A vssd1 vssd1 vccd1 vccd1 _5237_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5521_ _5524_/A _5539_/A vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__xor2_2
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5452_ _5454_/A _5454_/B _5451_/X vssd1 vssd1 vccd1 vccd1 _5576_/B sky130_fd_sc_hd__a21o_1
X_4403_ _4403_/A _4403_/B vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__xnor2_4
X_5383_ _5385_/A _5385_/B _5382_/Y vssd1 vssd1 vccd1 vccd1 _5384_/B sky130_fd_sc_hd__a21oi_2
X_4334_ _5486_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4335_/B sky130_fd_sc_hd__and3_2
XFILLER_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4265_ _4265_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__xor2_1
X_6004_ _6000_/B _6004_/B vssd1 vssd1 vccd1 vccd1 _6004_/X sky130_fd_sc_hd__and2b_1
X_4196_ _4223_/A _4223_/B _4195_/A vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__o21ai_1
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3216_ _3216_/A vssd1 vssd1 vccd1 vccd1 _3216_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _5720_/A _5720_/B vssd1 vssd1 vccd1 vccd1 _5719_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ _4050_/A _4472_/A vssd1 vssd1 vccd1 vccd1 _4474_/C sky130_fd_sc_hd__nand2_2
Xinput6 io_in[8] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4951_/A _4951_/B _4951_/C vssd1 vssd1 vccd1 vccd1 _5193_/B sky130_fd_sc_hd__a21oi_2
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ _5122_/A _3903_/B _3903_/C vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__and3_1
X_4883_ _4866_/B _4868_/X _4882_/A _4909_/A vssd1 vssd1 vccd1 vccd1 _4951_/B sky130_fd_sc_hd__o211ai_2
X_3834_ _5015_/A _3849_/B vssd1 vssd1 vccd1 vccd1 _3856_/A sky130_fd_sc_hd__and2_1
X_6622_ _6622_/A _3319_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_6553_ _6553_/A _3238_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
X_3765_ _3668_/B _3765_/B vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__and2b_1
X_3696_ _3696_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__xnor2_4
X_5504_ _5516_/A _5516_/B _5503_/Y vssd1 vssd1 vccd1 vccd1 _5506_/A sky130_fd_sc_hd__o21a_1
X_5435_ _5413_/X _5435_/B vssd1 vssd1 vccd1 vccd1 _5436_/B sky130_fd_sc_hd__and2b_1
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _5407_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5411_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4317_ _5428_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4318_/B sky130_fd_sc_hd__nand2_1
X_5297_ _5297_/A _5297_/B _5297_/C vssd1 vssd1 vccd1 vccd1 _5297_/X sky130_fd_sc_hd__and3_1
XFILLER_87_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4248_ _4251_/A _4251_/B vssd1 vssd1 vccd1 vccd1 _4248_/X sky130_fd_sc_hd__and2b_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4179_ _5350_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4180_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3550_ _3550_/A _3550_/B vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__or2_1
X_3481_ _3440_/B _3447_/A _3440_/A vssd1 vssd1 vccd1 vccd1 _3482_/B sky130_fd_sc_hd__o21ai_1
X_5220_ _5209_/Y _5217_/X _5218_/Y _5219_/X vssd1 vssd1 vccd1 vccd1 _5225_/A sky130_fd_sc_hd__a211oi_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5151_ _5151_/A _5151_/B vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__xnor2_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4102_ _4101_/A _4101_/B _4101_/C vssd1 vssd1 vccd1 vccd1 _4389_/C sky130_fd_sc_hd__a21o_1
X_5082_ _5147_/A _5147_/B _5081_/X vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4033_ _5353_/A vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _5984_/A vssd1 vssd1 vccd1 vccd1 _5997_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4935_ _4739_/A _4739_/B _4739_/C vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4866_ _4866_/A _4866_/B vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__nor2_2
X_3817_ _5356_/A _4174_/B _3810_/A vssd1 vssd1 vccd1 vccd1 _3817_/Y sky130_fd_sc_hd__a21boi_1
X_4797_ _4775_/A _4773_/Y _4769_/Y _4772_/X vssd1 vssd1 vccd1 vccd1 _4798_/B sky130_fd_sc_hd__o211a_1
X_6605_ _6605_/A _3300_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3748_ _4891_/B vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6536_ _6536_/A _3216_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
X_3679_ _4851_/A _3689_/B _3678_/X vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__o21a_2
X_5418_ _5419_/B _5418_/B vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__xnor2_2
X_6398_ _6401_/CLK _6398_/D vssd1 vssd1 vccd1 vccd1 _6398_/Q sky130_fd_sc_hd__dfxtp_1
X_5349_ _5458_/A _5322_/B _5255_/A _5322_/A vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__a22o_1
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4720_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4919_/B sky130_fd_sc_hd__xor2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4651_ _4651_/A _4891_/C vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__nand2_1
X_3602_ _3603_/A _3603_/B vssd1 vssd1 vccd1 vccd1 _3604_/A sky130_fd_sc_hd__nor2_1
X_4582_ _4905_/C _4600_/B _4580_/X _5711_/A _5712_/A vssd1 vssd1 vccd1 vccd1 _4583_/B
+ sky130_fd_sc_hd__o221a_1
X_3533_ _3718_/C vssd1 vssd1 vccd1 vccd1 _3716_/C sky130_fd_sc_hd__clkbuf_2
X_6321_ _6361_/CLK _6321_/D vssd1 vssd1 vccd1 vccd1 _6321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3464_ _3469_/B _3464_/B vssd1 vssd1 vccd1 vccd1 _3485_/B sky130_fd_sc_hd__nand2_1
X_6252_ _6256_/C _6294_/B vssd1 vssd1 vccd1 vccd1 _6402_/D sky130_fd_sc_hd__nor2_1
X_5203_ _5248_/A _5290_/B vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__nand2_1
X_6183_ _6375_/Q _6183_/B vssd1 vssd1 vccd1 vccd1 _6184_/A sky130_fd_sc_hd__and2_1
XFILLER_97_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3395_ _3395_/A _3395_/B _3430_/C vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__and3_1
X_5134_ _5134_/A _5134_/B vssd1 vssd1 vccd1 vccd1 _5135_/B sky130_fd_sc_hd__xor2_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5065_ _5065_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _5072_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4016_ _4016_/A _4016_/B vssd1 vssd1 vccd1 vccd1 _4016_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5967_ _5967_/A vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__clkbuf_2
X_4918_ _4792_/B _4918_/B vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5898_ _6423_/Q _5888_/Y _5892_/X _5893_/Y _5897_/Y vssd1 vssd1 vccd1 vccd1 _5898_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4849_ _4830_/B _4850_/B _4874_/C vssd1 vssd1 vccd1 vccd1 _4851_/B sky130_fd_sc_hd__a21o_1
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5821_ _5759_/Y _5818_/X _5820_/X _5758_/Y vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5752_ _5742_/A _5748_/X _5750_/X _5751_/Y vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__o22a_1
X_4703_ _4704_/A _4703_/B vssd1 vssd1 vccd1 vccd1 _4791_/B sky130_fd_sc_hd__xnor2_1
X_5683_ _5842_/A _5684_/B _5682_/X vssd1 vssd1 vccd1 vccd1 _5683_/X sky130_fd_sc_hd__a21o_1
X_4634_ _5743_/A vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4565_ _4565_/A _4565_/B vssd1 vssd1 vccd1 vccd1 _4565_/X sky130_fd_sc_hd__or2_1
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3516_ _3516_/A _3516_/B vssd1 vssd1 vccd1 vccd1 _3560_/B sky130_fd_sc_hd__xor2_1
X_6304_ _6304_/A _6309_/C vssd1 vssd1 vccd1 vccd1 _6304_/Y sky130_fd_sc_hd__nor2_1
X_4496_ _4496_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4497_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3447_ _3447_/A _3447_/B vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__or2_1
X_6235_ _6395_/Q _6243_/B vssd1 vssd1 vccd1 vccd1 _6236_/A sky130_fd_sc_hd__and2_1
X_3378_ _4711_/A vssd1 vssd1 vccd1 vccd1 _3395_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6183_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5117_ _5061_/A _5110_/A _5103_/Y _5105_/A vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__o22a_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6097_/A _6103_/C _6097_/C vssd1 vssd1 vccd1 vccd1 _6097_/X sky130_fd_sc_hd__and3_1
XFILLER_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5048_ _5048_/A _5048_/B vssd1 vssd1 vccd1 vccd1 _5049_/B sky130_fd_sc_hd__or2_1
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4354_/B sky130_fd_sc_hd__xnor2_1
X_3301_ _3303_/A vssd1 vssd1 vccd1 vccd1 _3301_/Y sky130_fd_sc_hd__inv_2
X_4281_ _4306_/A _4306_/B _4280_/A vssd1 vssd1 vccd1 vccd1 _4304_/B sky130_fd_sc_hd__o21bai_2
XFILLER_98_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3235_/A vssd1 vssd1 vccd1 vccd1 _3232_/Y sky130_fd_sc_hd__inv_2
X_6020_ _6001_/S _6017_/X _6018_/Y _4630_/A vssd1 vssd1 vccd1 vccd1 _6021_/B sky130_fd_sc_hd__a31o_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5804_ _5748_/B _5804_/B vssd1 vssd1 vccd1 vccd1 _5804_/X sky130_fd_sc_hd__and2b_1
X_3996_ _3996_/A _3996_/B _3996_/C vssd1 vssd1 vccd1 vccd1 _3996_/X sky130_fd_sc_hd__or3_4
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _5629_/Y _5634_/X _5645_/X _5733_/X _5734_/X vssd1 vssd1 vccd1 vccd1 _5774_/B
+ sky130_fd_sc_hd__a221o_1
X_5666_ _5666_/A _5666_/B _5666_/C vssd1 vssd1 vccd1 vccd1 _5671_/A sky130_fd_sc_hd__and3_1
X_4617_ _5789_/A _4617_/B _4617_/C _5789_/B vssd1 vssd1 vccd1 vccd1 _5805_/B sky130_fd_sc_hd__and4_2
X_5597_ _5596_/X _5595_/B _5593_/Y vssd1 vssd1 vccd1 vccd1 _5597_/Y sky130_fd_sc_hd__a21oi_1
X_4548_ _5684_/A _4550_/B _4547_/X vssd1 vssd1 vccd1 vccd1 _4549_/B sky130_fd_sc_hd__a21o_1
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4479_ _4487_/A _4487_/B _4478_/X vssd1 vssd1 vccd1 vccd1 _4479_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6218_ _6389_/Q _6232_/B vssd1 vssd1 vccd1 vccd1 _6219_/A sky130_fd_sc_hd__and2_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6149_ _6149_/A vssd1 vssd1 vccd1 vccd1 _6363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3850_ _3798_/B _3844_/A _3849_/Y vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__a21oi_1
X_3781_ _5371_/A vssd1 vssd1 vccd1 vccd1 _5316_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520_ _5538_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5539_/A sky130_fd_sc_hd__nand2_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5451_ _5450_/A _5451_/B vssd1 vssd1 vccd1 vccd1 _5451_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4402_ _4455_/A _4455_/B vssd1 vssd1 vccd1 vccd1 _4533_/A sky130_fd_sc_hd__xor2_4
X_5382_ _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5382_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4333_ _4333_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__nor2_2
X_4264_ _4288_/A _4288_/B vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__xor2_2
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3215_ _3216_/A vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__inv_2
X_6003_ _6003_/A vssd1 vssd1 vccd1 vccd1 _6330_/D sky130_fd_sc_hd__clkbuf_1
X_4195_ _4195_/A _4195_/B vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__nand2_1
XFILLER_94_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _3977_/A _3977_/B _4027_/A vssd1 vssd1 vccd1 vccd1 _3981_/C sky130_fd_sc_hd__a21bo_1
X_5718_ _5761_/A _5704_/B _5703_/A vssd1 vssd1 vccd1 vccd1 _5720_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _5622_/A _5622_/B _5228_/A vssd1 vssd1 vccd1 vccd1 _5650_/B sky130_fd_sc_hd__o21ai_2
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 io_in[9] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _4951_/A _4951_/B _4951_/C vssd1 vssd1 vccd1 vccd1 _5193_/A sky130_fd_sc_hd__and3_1
XFILLER_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3902_ _5154_/A _3931_/A vssd1 vssd1 vccd1 vccd1 _3903_/C sky130_fd_sc_hd__and2_1
XFILLER_60_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4882_ _4882_/A _4882_/B _4882_/C vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__nand3_2
X_6621_ _6621_/A _3318_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_3833_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3764_ _3961_/A _3961_/B _3763_/X vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__a21o_1
X_6552_ _6552_/A _3237_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
X_3695_ _3680_/Y _3697_/B _3694_/X vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__a21o_2
X_5503_ _5503_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _5503_/Y sky130_fd_sc_hd__nand2_1
X_5434_ _5434_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5465_/A sky130_fd_sc_hd__xnor2_2
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5365_ _5365_/A _5365_/B vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__nand2_1
X_4316_ _4327_/A _4327_/B vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5296_ _5296_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__nand2_1
X_4247_ _4247_/A _4247_/B vssd1 vssd1 vccd1 vccd1 _4251_/B sky130_fd_sc_hd__xnor2_2
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4178_ _4178_/A _4178_/B vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__xor2_1
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6485__67 vssd1 vssd1 vccd1 vccd1 _6485__67/HI _6593_/A sky130_fd_sc_hd__conb_1
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3480_ _3480_/A _3480_/B vssd1 vssd1 vccd1 vccd1 _3518_/A sky130_fd_sc_hd__xor2_2
X_5150_ _5150_/A _5596_/A vssd1 vssd1 vccd1 vccd1 _5654_/A sky130_fd_sc_hd__xnor2_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4101_ _4101_/A _4101_/B _4101_/C vssd1 vssd1 vccd1 vccd1 _4389_/B sky130_fd_sc_hd__nand3_2
X_5081_ _5076_/B _5081_/B vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__and2b_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4032_ _5560_/A vssd1 vssd1 vccd1 vccd1 _5353_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5983_ _5978_/A _5982_/A _5982_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _6327_/D sky130_fd_sc_hd__o211a_1
X_4934_ _4934_/A _4934_/B vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4865_ _4862_/X _4863_/X _4866_/A _4864_/Y vssd1 vssd1 vccd1 vccd1 _4866_/B sky130_fd_sc_hd__a211oi_2
X_6604_ _6604_/A _3299_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_3816_ _4152_/B vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__clkbuf_4
X_4796_ _4796_/A _4796_/B vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__xnor2_1
X_3747_ _3747_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _4131_/A sky130_fd_sc_hd__xor2_1
X_6535_ _6535_/A _3215_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_21_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3678_ _4828_/B _3677_/B vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__or2b_1
X_5417_ _5432_/A _5432_/B _5416_/X vssd1 vssd1 vccd1 vccd1 _5418_/B sky130_fd_sc_hd__a21oi_1
X_6397_ _6401_/CLK _6397_/D vssd1 vssd1 vccd1 vccd1 _6397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5348_ _5348_/A _5348_/B vssd1 vssd1 vccd1 vccd1 _5580_/B sky130_fd_sc_hd__xnor2_4
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5279_ _5535_/B vssd1 vssd1 vccd1 vccd1 _5458_/B sky130_fd_sc_hd__buf_2
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4650_ _4873_/B vssd1 vssd1 vccd1 vccd1 _4891_/C sky130_fd_sc_hd__clkbuf_2
X_3601_ _3605_/A _3605_/B _3600_/X vssd1 vssd1 vccd1 vccd1 _3603_/B sky130_fd_sc_hd__a21oi_1
X_4581_ _4581_/A vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__buf_4
X_6320_ _6361_/CLK _6320_/D vssd1 vssd1 vccd1 vccd1 _6320_/Q sky130_fd_sc_hd__dfxtp_1
X_3532_ _5815_/A _3409_/B _6038_/A vssd1 vssd1 vccd1 vccd1 _3718_/C sky130_fd_sc_hd__a21o_2
X_3463_ _3463_/A _3489_/A vssd1 vssd1 vccd1 vccd1 _3464_/B sky130_fd_sc_hd__nand2_1
X_6251_ _6402_/Q vssd1 vssd1 vccd1 vccd1 _6256_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5202_ _5297_/A _5202_/B vssd1 vssd1 vccd1 vccd1 _5205_/A sky130_fd_sc_hd__nand2_1
X_6182_ _6182_/A vssd1 vssd1 vccd1 vccd1 _6375_/D sky130_fd_sc_hd__clkbuf_1
X_5133_ _5126_/A _5126_/B _5132_/X vssd1 vssd1 vccd1 vccd1 _5145_/A sky130_fd_sc_hd__a21oi_2
X_3394_ _4763_/A _3592_/D vssd1 vssd1 vccd1 vccd1 _3430_/C sky130_fd_sc_hd__and2_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5064_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__nand2_1
X_4015_ _5237_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _6325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4917_ _4950_/A _4950_/B _4915_/Y _4916_/X vssd1 vssd1 vccd1 vccd1 _4948_/C sky130_fd_sc_hd__a211o_2
X_5897_ _5893_/Y _5892_/X _5896_/Y vssd1 vssd1 vccd1 vccd1 _5897_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4848_ _4831_/B _4842_/A _4831_/A vssd1 vssd1 vccd1 vccd1 _4852_/B sky130_fd_sc_hd__a21oi_1
X_4779_ _4779_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4779_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6455__37 vssd1 vssd1 vccd1 vccd1 _6455__37/HI _6560_/A sky130_fd_sc_hd__conb_1
XFILLER_113_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5820_ _5868_/C vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5751_ _5871_/B _5817_/A _5871_/A vssd1 vssd1 vccd1 vccd1 _5751_/Y sky130_fd_sc_hd__o21ai_2
X_4702_ _4706_/B _4702_/B vssd1 vssd1 vccd1 vccd1 _4703_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5682_ _5681_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5682_/X sky130_fd_sc_hd__and2b_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _5868_/A vssd1 vssd1 vccd1 vccd1 _5743_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4564_ _4562_/A _4562_/B _4563_/Y vssd1 vssd1 vccd1 vccd1 _4565_/B sky130_fd_sc_hd__o21ai_1
X_3515_ _3515_/A _3515_/B vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__nor2_1
X_6303_ _6422_/Q _6421_/Q _6303_/C vssd1 vssd1 vccd1 vccd1 _6309_/C sky130_fd_sc_hd__and3_1
XFILLER_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4495_ _4472_/X _4495_/B vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__and2b_1
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6234_ _6234_/A vssd1 vssd1 vccd1 vccd1 _6243_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3446_ _4924_/A _3509_/B _3446_/C vssd1 vssd1 vccd1 vccd1 _3447_/B sky130_fd_sc_hd__and3_1
X_3377_ _4677_/A vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/A vssd1 vssd1 vccd1 vccd1 _6369_/D sky130_fd_sc_hd__clkbuf_1
X_5116_ _5174_/A _5174_/B _5115_/X vssd1 vssd1 vccd1 vccd1 _5127_/A sky130_fd_sc_hd__o21bai_2
XFILLER_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6103_/A _6103_/B vssd1 vssd1 vccd1 vccd1 _6097_/C sky130_fd_sc_hd__xnor2_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5047_ _5048_/A _5048_/B vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5949_ _5945_/A _5909_/X _5946_/Y _5947_/X _5948_/X vssd1 vssd1 vccd1 vccd1 _6321_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3300_ _3303_/A vssd1 vssd1 vccd1 vccd1 _3300_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4280_ _4280_/A _4280_/B vssd1 vssd1 vccd1 vccd1 _4306_/B sky130_fd_sc_hd__or2_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3231_ _3235_/A vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__inv_2
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5803_ _5803_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__nand2_1
X_3995_ _3981_/A _3981_/B _3981_/C vssd1 vssd1 vccd1 vccd1 _3996_/C sky130_fd_sc_hd__a21oi_1
X_5734_ _5633_/A _5633_/B _5644_/Y _5637_/X vssd1 vssd1 vccd1 vccd1 _5734_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5665_ _5666_/A _5666_/B _5666_/C vssd1 vssd1 vccd1 vccd1 _5665_/X sky130_fd_sc_hd__a21o_1
X_4616_ _4506_/Y _5776_/A _5776_/B _5778_/A _4615_/Y vssd1 vssd1 vccd1 vccd1 _5789_/B
+ sky130_fd_sc_hd__o311a_2
X_5596_ _5596_/A _5150_/A vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__or2b_1
XFILLER_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ _4547_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4547_/X sky130_fd_sc_hd__and2_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4478_ _4003_/A _4003_/B _4004_/A vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__o21a_1
X_3429_ _4800_/A vssd1 vssd1 vccd1 vccd1 _4886_/A sky130_fd_sc_hd__buf_2
X_6217_ _6217_/A vssd1 vssd1 vccd1 vccd1 _6389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6148_ _6362_/Q _6164_/B vssd1 vssd1 vccd1 vccd1 _6149_/A sky130_fd_sc_hd__and2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6079_ _6078_/B _6078_/C _6078_/A vssd1 vssd1 vccd1 vccd1 _6083_/B sky130_fd_sc_hd__o21ai_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _5441_/A vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__clkbuf_2
X_5450_ _5450_/A _5451_/B vssd1 vssd1 vccd1 vccd1 _5454_/B sky130_fd_sc_hd__xnor2_2
X_4401_ _4399_/A _4399_/B _4400_/X vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__o21a_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5381_ _5382_/A _5382_/B vssd1 vssd1 vccd1 vccd1 _5385_/B sky130_fd_sc_hd__xor2_4
X_4332_ _5487_/A _4332_/B _4332_/C vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__and3_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6345_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_115_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4263_ _5560_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4288_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3214_ _3216_/A vssd1 vssd1 vccd1 vccd1 _3214_/Y sky130_fd_sc_hd__inv_2
X_6002_ _6134_/A _6002_/B vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__and2_1
X_4194_ _4194_/A _4194_/B vssd1 vssd1 vccd1 vccd1 _4195_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3978_ _3978_/A _3978_/B _3978_/C vssd1 vssd1 vccd1 vccd1 _4027_/A sky130_fd_sc_hd__nand3_1
XFILLER_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5717_ _5785_/A _5717_/B vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5648_ _5648_/A _5648_/B vssd1 vssd1 vccd1 vccd1 _5650_/A sky130_fd_sc_hd__nand2_2
X_5579_ _5640_/A _5640_/B _5578_/X vssd1 vssd1 vccd1 vccd1 _5636_/B sky130_fd_sc_hd__a21o_1
XFILLER_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4950_ _4950_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _5106_/A sky130_fd_sc_hd__xor2_4
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3901_ _5017_/A _4174_/B _3937_/B _3900_/A vssd1 vssd1 vccd1 vccd1 _3917_/B sky130_fd_sc_hd__a31o_1
X_4881_ _4878_/A _4878_/B _4878_/C vssd1 vssd1 vccd1 vccd1 _4882_/C sky130_fd_sc_hd__a21o_1
X_6620_ _6620_/A _3317_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_3832_ _5118_/A vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6551_ _6551_/A _3235_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_3763_ _3696_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__and2b_1
X_5502_ _5503_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _5516_/B sky130_fd_sc_hd__xnor2_2
X_3694_ _3693_/B _3694_/B vssd1 vssd1 vccd1 vccd1 _3694_/X sky130_fd_sc_hd__and2b_1
X_5433_ _5433_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5434_/B sky130_fd_sc_hd__nand2_1
X_5364_ _5364_/A _5364_/B vssd1 vssd1 vccd1 vccd1 _5365_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4315_ _4329_/A _4329_/B _4313_/A vssd1 vssd1 vccd1 vccd1 _4327_/B sky130_fd_sc_hd__o21a_1
XFILLER_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5295_ _5295_/A _5295_/B vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__xnor2_2
X_4246_ _4246_/A _4246_/B vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__xor2_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4177_ _4177_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4100_ _4100_/A _4100_/B vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5592_/A _5080_/B vssd1 vssd1 vccd1 vccd1 _5147_/B sky130_fd_sc_hd__and2_1
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4031_ _5555_/C vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5982_ _5982_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5982_/Y sky130_fd_sc_hd__nand2_1
X_4933_ _4941_/B vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__clkinv_2
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4864_ _4861_/A _4861_/C _4861_/B vssd1 vssd1 vccd1 vccd1 _4864_/Y sky130_fd_sc_hd__a21oi_1
X_3815_ _3960_/A _4152_/B vssd1 vssd1 vccd1 vccd1 _3875_/A sky130_fd_sc_hd__nand2_2
X_4795_ _4793_/X _4795_/B vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__and2b_1
X_6603_ _6603_/A _3297_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_3746_ _3757_/A _3757_/B _3757_/C vssd1 vssd1 vccd1 vccd1 _4101_/B sky130_fd_sc_hd__a21o_1
X_6534_ _6534_/A _3214_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5416_ _5415_/B _5416_/B vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__and2b_1
X_3677_ _4828_/B _3677_/B vssd1 vssd1 vccd1 vccd1 _3689_/B sky130_fd_sc_hd__xor2_1
X_6396_ _6396_/CLK _6396_/D vssd1 vssd1 vccd1 vccd1 _6396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5347_ _5583_/A _5583_/B vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__xor2_4
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5278_ _5424_/B vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4229_ _4404_/A _4957_/C _4184_/A _4228_/X vssd1 vssd1 vccd1 vccd1 _4383_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3600_ _3599_/B _3600_/B vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__and2b_1
X_4580_ _4596_/C _4580_/B vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__xor2_1
X_3531_ _6337_/Q vssd1 vssd1 vccd1 vccd1 _6038_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3462_ _3462_/A _3473_/C vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__and2_1
X_6250_ _6394_/Q _6395_/Q _6100_/X _6246_/X _6249_/X vssd1 vssd1 vccd1 vccd1 _6401_/D
+ sky130_fd_sc_hd__a41o_1
X_5201_ _5201_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__xnor2_1
X_6181_ _6228_/A input2/X vssd1 vssd1 vccd1 vccd1 _6182_/A sky130_fd_sc_hd__and2_1
X_3393_ _4642_/D vssd1 vssd1 vccd1 vccd1 _3592_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_111_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5132_ _5120_/A _5132_/B vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__and2b_1
XFILLER_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5063_ _5017_/A _5297_/B _5001_/A _5062_/X vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__a31o_1
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4014_ _4014_/A _4109_/B vssd1 vssd1 vccd1 vccd1 _4014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5965_ _6365_/Q _6025_/B vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__and2_1
X_4916_ _4846_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__and2b_1
X_5896_ _6425_/Q _5896_/B vssd1 vssd1 vccd1 vccd1 _5896_/Y sky130_fd_sc_hd__nor2_1
X_4847_ _4847_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4913_/B sky130_fd_sc_hd__xnor2_4
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4778_ _4789_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__xor2_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3729_ _3729_/A _3735_/B vssd1 vssd1 vccd1 vccd1 _3731_/B sky130_fd_sc_hd__nand2_1
X_6379_ _6388_/CLK _6379_/D vssd1 vssd1 vccd1 vccd1 _6379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6522__104 vssd1 vssd1 vccd1 vccd1 _6522__104/HI _6630_/A sky130_fd_sc_hd__conb_1
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5750_ _5750_/A _5750_/B vssd1 vssd1 vccd1 vccd1 _5750_/X sky130_fd_sc_hd__xor2_2
X_4701_ _4701_/A _4701_/B vssd1 vssd1 vccd1 vccd1 _4702_/B sky130_fd_sc_hd__xnor2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5681_/A _5682_/B vssd1 vssd1 vccd1 vccd1 _5684_/B sky130_fd_sc_hd__xnor2_1
X_4632_ _5745_/A vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _5785_/A _4586_/B vssd1 vssd1 vccd1 vccd1 _4563_/Y sky130_fd_sc_hd__nand2_1
X_3514_ _3516_/A _3516_/B vssd1 vssd1 vccd1 vccd1 _3518_/B sky130_fd_sc_hd__or2b_1
X_6302_ _6421_/Q _6303_/C _6301_/Y vssd1 vssd1 vccd1 vccd1 _6421_/D sky130_fd_sc_hd__o21a_1
X_4494_ _5790_/A vssd1 vssd1 vccd1 vccd1 _4617_/C sky130_fd_sc_hd__inv_2
X_3445_ _3445_/A _3445_/B vssd1 vssd1 vccd1 vccd1 _3791_/A sky130_fd_sc_hd__or2_2
X_6233_ _6233_/A vssd1 vssd1 vccd1 vccd1 _6395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3376_ _4745_/A vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6368_/Q _6164_/B vssd1 vssd1 vccd1 vccd1 _6165_/A sky130_fd_sc_hd__and2_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5115_ _5112_/A _5115_/B vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__and2b_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6095_ _6104_/B _6032_/X _6094_/X _5948_/X vssd1 vssd1 vccd1 vccd1 _6344_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5046_ _5046_/A vssd1 vssd1 vccd1 vccd1 _5048_/B sky130_fd_sc_hd__inv_2
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5948_ _6115_/B vssd1 vssd1 vccd1 vccd1 _5948_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5879_ _6418_/Q vssd1 vssd1 vccd1 vccd1 _6294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6515__97 vssd1 vssd1 vccd1 vccd1 _6515__97/HI _6623_/A sky130_fd_sc_hd__conb_1
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6427__9 vssd1 vssd1 vccd1 vccd1 _6427__9/HI _6532_/A sky130_fd_sc_hd__conb_1
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3230_ _3248_/A vssd1 vssd1 vccd1 vccd1 _3235_/A sky130_fd_sc_hd__buf_12
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5802_ _5784_/X _5794_/X _5801_/X vssd1 vssd1 vccd1 vccd1 _5802_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3994_ _4005_/A _3994_/B vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__or2_1
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5733_ _5659_/X _5670_/X _5729_/X _5730_/Y _5732_/X vssd1 vssd1 vccd1 vccd1 _5733_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5664_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5666_/C sky130_fd_sc_hd__xnor2_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4615_ _5769_/A vssd1 vssd1 vccd1 vccd1 _4615_/Y sky130_fd_sc_hd__inv_2
X_5595_ _5593_/Y _5595_/B vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__and2b_2
X_4546_ _4547_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4550_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4477_ _4487_/A _4487_/B _4476_/X vssd1 vssd1 vccd1 vccd1 _4488_/B sky130_fd_sc_hd__o21bai_1
X_3428_ _3646_/A vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__clkbuf_2
X_6216_ _6388_/Q _6232_/B vssd1 vssd1 vccd1 vccd1 _6217_/A sky130_fd_sc_hd__and2_1
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6147_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6164_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3359_ _3359_/A vssd1 vssd1 vccd1 vccd1 _3409_/B sky130_fd_sc_hd__buf_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6078_ _6078_/A _6078_/B _6078_/C vssd1 vssd1 vccd1 vccd1 _6078_/X sky130_fd_sc_hd__or3_1
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5029_ _5937_/A _5029_/B _5029_/C vssd1 vssd1 vccd1 vccd1 _5035_/B sky130_fd_sc_hd__and3_1
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _4403_/A _4403_/B vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__or2b_1
X_5380_ _5398_/A _5398_/B _5379_/X vssd1 vssd1 vccd1 vccd1 _5382_/B sky130_fd_sc_hd__a21oi_2
X_4331_ _5487_/A _4332_/B _4332_/C vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__a21oi_1
X_4262_ _4262_/A _4262_/B vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__xnor2_2
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3213_ _3216_/A vssd1 vssd1 vccd1 vccd1 _3213_/Y sky130_fd_sc_hd__clkinv_4
X_6001_ _4629_/B _6000_/Y _6001_/S vssd1 vssd1 vccd1 vccd1 _6002_/B sky130_fd_sc_hd__mux2_1
X_6528__110 vssd1 vssd1 vccd1 vccd1 _6528__110/HI _6636_/A sky130_fd_sc_hd__conb_1
X_4193_ _4194_/A _4194_/B vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__or2_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3977_ _3977_/A _3977_/B vssd1 vssd1 vccd1 vccd1 _3978_/C sky130_fd_sc_hd__xor2_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5716_ _5704_/Y _5714_/Y _5715_/Y vssd1 vssd1 vccd1 vccd1 _5716_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5647_ _5647_/A vssd1 vssd1 vccd1 vccd1 _5648_/B sky130_fd_sc_hd__inv_2
X_5578_ _5421_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4529_ _5790_/A _4562_/A vssd1 vssd1 vccd1 vccd1 _4529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3900_ _3900_/A _3900_/B vssd1 vssd1 vccd1 vccd1 _3937_/B sky130_fd_sc_hd__nor2_1
X_4880_ _4624_/A _4891_/C _4875_/B _4879_/Y vssd1 vssd1 vccd1 vccd1 _4882_/B sky130_fd_sc_hd__a31o_1
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3831_ _5154_/A vssd1 vssd1 vccd1 vccd1 _5118_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6550_ _6550_/A _3234_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_3762_ _4010_/A _4010_/B _3761_/Y vssd1 vssd1 vccd1 vccd1 _3961_/B sky130_fd_sc_hd__a21bo_2
XFILLER_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5501_ _5517_/A _5517_/B vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__and2_1
X_3693_ _3694_/B _3693_/B vssd1 vssd1 vccd1 vccd1 _3697_/B sky130_fd_sc_hd__xnor2_2
X_5432_ _5432_/A _5432_/B vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__xnor2_2
X_5363_ _5363_/A _5363_/B vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__xor2_2
X_4314_ _4314_/A _4314_/B vssd1 vssd1 vccd1 vccd1 _4329_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5294_ _5294_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5295_/B sky130_fd_sc_hd__xnor2_2
X_4245_ _4218_/A _4218_/B _4244_/Y vssd1 vssd1 vccd1 vccd1 _4251_/A sky130_fd_sc_hd__o21ba_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4176_ _4581_/A _3958_/B _4173_/A _4200_/A vssd1 vssd1 vccd1 vccd1 _4207_/A sky130_fd_sc_hd__a31oi_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6476__58 vssd1 vssd1 vccd1 vccd1 _6476__58/HI _6584_/A sky130_fd_sc_hd__conb_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4030_ _4373_/A vssd1 vssd1 vccd1 vccd1 _5555_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _5981_/A _5981_/B vssd1 vssd1 vccd1 vccd1 _5982_/B sky130_fd_sc_hd__xnor2_1
X_4932_ _4981_/S _4932_/B vssd1 vssd1 vccd1 vccd1 _4941_/B sky130_fd_sc_hd__and2_1
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6602_ _6602_/A _3341_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_4863_ _4863_/A _4857_/B vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__or2b_1
X_3814_ _4021_/B vssd1 vssd1 vccd1 vccd1 _4152_/B sky130_fd_sc_hd__clkbuf_2
X_4794_ _4794_/A _4794_/B _4794_/C vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__or3_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6533_ _6533_/A _3213_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
X_3745_ _3747_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3757_/C sky130_fd_sc_hd__nand2_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5415_ _5416_/B _5415_/B vssd1 vssd1 vccd1 vccd1 _5432_/B sky130_fd_sc_hd__xnor2_2
X_3676_ _3683_/B _3703_/B _3683_/A vssd1 vssd1 vccd1 vccd1 _3677_/B sky130_fd_sc_hd__a21bo_1
X_6395_ _6396_/CLK _6395_/D vssd1 vssd1 vccd1 vccd1 _6395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _5346_/A _5346_/B vssd1 vssd1 vccd1 vccd1 _5583_/B sky130_fd_sc_hd__and2_1
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5277_ _5275_/Y _5276_/X _5231_/C vssd1 vssd1 vccd1 vccd1 _5424_/B sky130_fd_sc_hd__a21oi_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4228_ _4624_/A _4957_/B _3589_/A vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__or3b_1
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4159_ _4150_/X _4157_/X _4121_/Y _4158_/X vssd1 vssd1 vccd1 vccd1 _4159_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6490__72 vssd1 vssd1 vccd1 vccd1 _6490__72/HI _6598_/A sky130_fd_sc_hd__conb_1
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3530_ _4850_/A vssd1 vssd1 vccd1 vccd1 _4888_/A sky130_fd_sc_hd__buf_2
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3461_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3473_/C sky130_fd_sc_hd__inv_2
X_5200_ _5201_/B _5201_/A vssd1 vssd1 vccd1 vccd1 _5207_/A sky130_fd_sc_hd__and2b_1
X_6180_ _6100_/X _6175_/X _6176_/X _6179_/X vssd1 vssd1 vccd1 vccd1 _6374_/D sky130_fd_sc_hd__a31o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3392_ _3356_/A _6345_/Q _6341_/Q vssd1 vssd1 vccd1 vccd1 _4642_/D sky130_fd_sc_hd__a21o_1
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _5127_/A _5127_/B _5153_/A vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__a21bo_1
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5062_ _5064_/A _5299_/B _5119_/B vssd1 vssd1 vccd1 vccd1 _5062_/X sky130_fd_sc_hd__and3_1
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4013_ _4373_/B vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5964_ _5964_/A vssd1 vssd1 vccd1 vccd1 _6324_/D sky130_fd_sc_hd__clkbuf_1
X_4915_ _4824_/B _4824_/C _4824_/A vssd1 vssd1 vccd1 vccd1 _4915_/Y sky130_fd_sc_hd__a21oi_1
X_5895_ _3354_/X _5870_/X _5894_/X _4634_/X vssd1 vssd1 vccd1 vccd1 _5896_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _4846_/A _4916_/B vssd1 vssd1 vccd1 vccd1 _4950_/A sky130_fd_sc_hd__xnor2_4
X_4777_ _4777_/A _4777_/B vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__xor2_1
X_3728_ _3730_/A _3730_/C _3736_/A vssd1 vssd1 vccd1 vccd1 _3732_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3659_ _6327_/Q _3592_/C _4694_/B _6326_/Q vssd1 vssd1 vccd1 vccd1 _3660_/B sky130_fd_sc_hd__a22oi_1
X_6378_ _6388_/CLK _6378_/D vssd1 vssd1 vccd1 vccd1 _6378_/Q sky130_fd_sc_hd__dfxtp_1
X_5329_ _5326_/A _5326_/B _5327_/B _5328_/Y vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__a31o_2
XFILLER_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6446__28 vssd1 vssd1 vccd1 vccd1 _6446__28/HI _6551_/A sky130_fd_sc_hd__conb_1
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4700_ _4700_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4701_/B sky130_fd_sc_hd__xor2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5680_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4631_ _5756_/A _5979_/A _5756_/C _5756_/D vssd1 vssd1 vccd1 vccd1 _5745_/A sky130_fd_sc_hd__nor4_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4562_ _4562_/A _4562_/B vssd1 vssd1 vccd1 vccd1 _4586_/B sky130_fd_sc_hd__xor2_1
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3513_ _3513_/A _3520_/A vssd1 vssd1 vccd1 vccd1 _3516_/B sky130_fd_sc_hd__nand2_1
X_4493_ _4493_/A _4493_/B vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__xnor2_4
X_6301_ _6304_/A _6301_/B vssd1 vssd1 vccd1 vccd1 _6301_/Y sky130_fd_sc_hd__nor2_1
X_3444_ _3482_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3445_/B sky130_fd_sc_hd__nor2_1
X_6232_ _6394_/Q _6232_/B vssd1 vssd1 vccd1 vccd1 _6233_/A sky130_fd_sc_hd__and2_1
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6163_/A vssd1 vssd1 vccd1 vccd1 _6368_/D sky130_fd_sc_hd__clkbuf_1
X_3375_ _6333_/Q vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5114_ _5114_/A _5114_/B vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__xor2_2
XFILLER_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6092_/X _6103_/C _6036_/A vssd1 vssd1 vccd1 vccd1 _6094_/X sky130_fd_sc_hd__a21bo_1
XFILLER_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A _5045_/B vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6460__42 vssd1 vssd1 vccd1 vccd1 _6460__42/HI _6565_/A sky130_fd_sc_hd__conb_1
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _5946_/A _5946_/B _5933_/B vssd1 vssd1 vccd1 vccd1 _5947_/X sky130_fd_sc_hd__a21bo_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5878_ _6419_/Q _6418_/Q _5875_/X _5877_/Y vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__o31a_1
X_4829_ _4830_/B _4830_/C _4830_/D _4830_/A vssd1 vssd1 vccd1 vccd1 _4831_/B sky130_fd_sc_hd__a22o_1
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _6405_/Q _5792_/X _5800_/X _6406_/Q vssd1 vssd1 vccd1 vccd1 _5801_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3993_ _4581_/A _4041_/B _3992_/C vssd1 vssd1 vccd1 vccd1 _3994_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5732_ _5731_/A _5657_/Y _5659_/A _5731_/X vssd1 vssd1 vccd1 vccd1 _5732_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5663_ _5663_/A _5529_/Y vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__or2b_1
X_4614_ _4614_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__or2_2
X_5594_ _5593_/A _5593_/B _5593_/C vssd1 vssd1 vccd1 vccd1 _5595_/B sky130_fd_sc_hd__o21ai_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4545_ _4545_/A _4545_/B vssd1 vssd1 vccd1 vccd1 _4547_/B sky130_fd_sc_hd__and2_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4476_ _4476_/A _4476_/B vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__xor2_1
X_6215_ _6234_/A vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3427_ _6329_/Q vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6146_ _6146_/A vssd1 vssd1 vccd1 vccd1 _6362_/D sky130_fd_sc_hd__clkbuf_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _6345_/Q vssd1 vssd1 vccd1 vccd1 _3359_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3289_ _3291_/A vssd1 vssd1 vccd1 vccd1 _3289_/Y sky130_fd_sc_hd__inv_2
X_6077_ _6063_/Y _6077_/B vssd1 vssd1 vccd1 vccd1 _6078_/C sky130_fd_sc_hd__and2b_1
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5028_/A _5040_/B _5031_/A vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__and3_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _4383_/A _4330_/B vssd1 vssd1 vccd1 vccd1 _4332_/C sky130_fd_sc_hd__and2_1
XFILLER_5_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ _5362_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4262_/B sky130_fd_sc_hd__nand2_1
X_3212_ _3216_/A vssd1 vssd1 vccd1 vccd1 _3212_/Y sky130_fd_sc_hd__inv_2
X_6000_ _6004_/B _6000_/B vssd1 vssd1 vccd1 vccd1 _6000_/Y sky130_fd_sc_hd__xnor2_1
X_4192_ _4014_/A _4183_/X _4188_/X _4225_/A vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__a31oi_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6430__12 vssd1 vssd1 vccd1 vccd1 _6430__12/HI _6535_/A sky130_fd_sc_hd__conb_1
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3976_ _3975_/A _3991_/A _5068_/A _4118_/B vssd1 vssd1 vccd1 vccd1 _3978_/B sky130_fd_sc_hd__a2bb2o_1
X_5715_ _5916_/A _5710_/Y _5714_/B _5714_/A vssd1 vssd1 vccd1 vccd1 _5715_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5646_ _5738_/A _5695_/A vssd1 vssd1 vccd1 vccd1 _5659_/A sky130_fd_sc_hd__xor2_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5577_ _5655_/A _5655_/B _5576_/X vssd1 vssd1 vccd1 vccd1 _5640_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4528_ _5759_/A _4569_/A vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__or2_1
X_4459_ _4353_/B _4459_/B vssd1 vssd1 vccd1 vccd1 _4459_/X sky130_fd_sc_hd__and2b_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6129_ _6347_/Q _6350_/Q _6129_/C vssd1 vssd1 vccd1 vccd1 _6129_/X sky130_fd_sc_hd__and3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _5198_/A vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__clkbuf_2
X_3761_ _3761_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3761_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5500_ _5500_/A _5500_/B vssd1 vssd1 vccd1 vccd1 _5517_/B sky130_fd_sc_hd__nor2_2
X_3692_ _3692_/A _3707_/A vssd1 vssd1 vccd1 vccd1 _3693_/B sky130_fd_sc_hd__and2_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5431_ _5296_/A _5560_/B _5434_/A _5430_/A vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__a31o_2
X_5362_ _5362_/A _5428_/B vssd1 vssd1 vccd1 vccd1 _5363_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4313_ _4313_/A _4313_/B vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5293_ _5330_/A _5330_/B _5292_/X vssd1 vssd1 vccd1 vccd1 _5295_/A sky130_fd_sc_hd__a21oi_2
XFILLER_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4244_ _4244_/A _4244_/B vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__nor2_1
X_4175_ _4208_/A _4208_/B vssd1 vssd1 vccd1 vccd1 _4200_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3959_ _3959_/A _3959_/B vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5629_ _5629_/A vssd1 vssd1 vccd1 vccd1 _5629_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5980_ _5978_/X _5980_/B vssd1 vssd1 vccd1 vccd1 _5981_/B sky130_fd_sc_hd__and2b_1
X_4931_ _4931_/A _4931_/B _4931_/C vssd1 vssd1 vccd1 vccd1 _4932_/B sky130_fd_sc_hd__or3_1
X_4862_ _4862_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__or2b_1
X_6601_ _6601_/A _3296_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_3813_ _3813_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__xor2_4
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4793_ _4794_/B _4794_/C _4794_/A vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3744_ _4682_/A _4957_/C _3754_/A _3743_/Y vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__o22ai_2
X_6532_ _6532_/A _3212_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
X_3675_ _6327_/Q _3646_/C _3699_/D _3672_/A vssd1 vssd1 vccd1 vccd1 _3683_/A sky130_fd_sc_hd__a22o_1
X_5414_ _5436_/A _5435_/B _5413_/X vssd1 vssd1 vccd1 vccd1 _5415_/B sky130_fd_sc_hd__a21oi_2
X_6394_ _6396_/CLK _6394_/D vssd1 vssd1 vccd1 vccd1 _6394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5345_ _5348_/A _5348_/B vssd1 vssd1 vccd1 vccd1 _5346_/B sky130_fd_sc_hd__or2b_1
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5276_ _5275_/B _4960_/A _4960_/B vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4227_ _4905_/A vssd1 vssd1 vccd1 vccd1 _4624_/A sky130_fd_sc_hd__clkbuf_2
X_4158_ _4121_/B _4121_/C _4121_/D _4121_/A vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4089_ _4089_/A _4470_/A vssd1 vssd1 vccd1 vccd1 _4472_/C sky130_fd_sc_hd__or2_1
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3460_ _4697_/A _4651_/A _3494_/B _3466_/B vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__and4_1
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3391_ _3653_/A vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5152_/A _5152_/B vssd1 vssd1 vccd1 vccd1 _5153_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5061_ _5061_/A _5061_/B vssd1 vssd1 vccd1 vccd1 _5119_/B sky130_fd_sc_hd__xor2_2
XFILLER_96_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4012_ _4340_/B vssd1 vssd1 vccd1 vccd1 _4373_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5963_ _6374_/Q _6025_/B vssd1 vssd1 vccd1 vccd1 _5964_/A sky130_fd_sc_hd__and2_1
X_4914_ _4963_/A _4963_/B _4913_/X vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__a21o_2
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5894_ _4619_/X _5823_/C _3364_/B _5742_/B vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__o2bb2a_1
X_4845_ _4845_/A _4844_/X vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__or2b_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4776_ _4776_/A _4768_/A vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__or2b_1
X_3727_ _3735_/A _3735_/B _3735_/C vssd1 vssd1 vccd1 vccd1 _3736_/A sky130_fd_sc_hd__a21oi_2
X_3658_ _3649_/A _3648_/B _3648_/C vssd1 vssd1 vccd1 vccd1 _3682_/B sky130_fd_sc_hd__a21o_1
X_3589_ _3589_/A _3589_/B vssd1 vssd1 vccd1 vccd1 _3589_/Y sky130_fd_sc_hd__nand2_1
X_6377_ _6396_/CLK _6377_/D vssd1 vssd1 vccd1 vccd1 _6377_/Q sky130_fd_sc_hd__dfxtp_1
X_5328_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5328_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5259_ _5296_/A _5350_/B _5259_/C vssd1 vssd1 vccd1 vccd1 _5267_/B sky130_fd_sc_hd__nand3_1
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4630_ _4630_/A _5967_/A _4630_/C vssd1 vssd1 vccd1 vccd1 _5756_/D sky130_fd_sc_hd__or3_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6300_ _6421_/Q _6303_/C vssd1 vssd1 vccd1 vccd1 _6301_/B sky130_fd_sc_hd__and2_1
X_4561_ _5067_/A vssd1 vssd1 vccd1 vccd1 _5785_/A sky130_fd_sc_hd__buf_2
X_3512_ _3519_/A _3519_/B vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__or2_1
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ _4476_/X _4479_/Y _4488_/B _4478_/X vssd1 vssd1 vccd1 vccd1 _4493_/B sky130_fd_sc_hd__o2bb2a_1
X_3443_ _3482_/A _3444_/B vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__and2_1
X_6231_ _6231_/A vssd1 vssd1 vccd1 vccd1 _6394_/D sky130_fd_sc_hd__clkbuf_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6367_/Q _6164_/B vssd1 vssd1 vccd1 vccd1 _6163_/A sky130_fd_sc_hd__and2_1
X_5113_ _5168_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3374_ _5017_/A vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6093_/A _6092_/A vssd1 vssd1 vccd1 vccd1 _6103_/C sky130_fd_sc_hd__or2b_1
XFILLER_84_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5946_ _5946_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5877_ _5765_/X _5870_/A _5876_/X _5807_/A vssd1 vssd1 vccd1 vccd1 _5877_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4828_ _4828_/A _4828_/B vssd1 vssd1 vccd1 vccd1 _4831_/A sky130_fd_sc_hd__xnor2_1
X_4759_ _4809_/A vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__inv_2
XFILLER_108_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6506__88 vssd1 vssd1 vccd1 vccd1 _6506__88/HI _6614_/A sky130_fd_sc_hd__conb_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3992_ _4581_/A _3992_/B _3992_/C vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__and3_1
X_5800_ _5936_/A _5746_/X _5799_/X _5743_/A vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__o2bb2a_1
X_5731_ _5731_/A _5731_/B vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__and2_1
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5662_ _5736_/B _5662_/B vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__xnor2_1
X_5593_ _5593_/A _5593_/B _5593_/C vssd1 vssd1 vccd1 vccd1 _5593_/Y sky130_fd_sc_hd__nor3_1
X_4613_ _5777_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__nand2_1
X_4544_ _4544_/A _4544_/B _4553_/A vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__or3_1
X_4475_ _4594_/B _4594_/C _4594_/A vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__a21boi_4
X_6214_ _6214_/A vssd1 vssd1 vccd1 vccd1 _6388_/D sky130_fd_sc_hd__clkbuf_1
X_3426_ _3426_/A _3426_/B vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__nor2_1
X_6145_ _6361_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6146_/A sky130_fd_sc_hd__and2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3409_/A vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__buf_2
X_6076_ _6341_/Q _6060_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__o21a_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5020_/B _5027_/B vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__and2b_1
X_3288_ _3291_/A vssd1 vssd1 vccd1 vccd1 _3288_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5929_ _6134_/A _5929_/B vssd1 vssd1 vccd1 vccd1 _5930_/A sky130_fd_sc_hd__and2_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _4212_/Y _4297_/A _4266_/A _4266_/B vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__o22a_1
XFILLER_113_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4191_ _5406_/A _4298_/B _4191_/C vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__and3_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3211_ _3342_/A vssd1 vssd1 vccd1 vccd1 _3216_/A sky130_fd_sc_hd__buf_6
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _3975_/A _3991_/A _5095_/A _4118_/B vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__or4bb_1
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5714_ _5714_/A _5714_/B vssd1 vssd1 vccd1 vccd1 _5714_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5645_ _5637_/X _5643_/Y _5644_/Y vssd1 vssd1 vccd1 vccd1 _5645_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5576_ _5453_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _5576_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4527_ _4527_/A _4527_/B vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__xnor2_4
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4458_ _4379_/X _4579_/B _4578_/A vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__a21o_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6497__79 vssd1 vssd1 vccd1 vccd1 _6497__79/HI _6605_/A sky130_fd_sc_hd__conb_1
X_3409_ _3409_/A _3409_/B vssd1 vssd1 vccd1 vccd1 _3472_/B sky130_fd_sc_hd__and2_1
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4389_ _5545_/A _4389_/B _4389_/C vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__and3_1
X_6128_ _6351_/Q _6352_/Q _6354_/Q _6353_/Q vssd1 vssd1 vccd1 vccd1 _6129_/C sky130_fd_sc_hd__and4_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6059_ _6059_/A vssd1 vssd1 vccd1 vccd1 _6074_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _3733_/X _3758_/X _4057_/A vssd1 vssd1 vccd1 vccd1 _4010_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3691_ _3692_/A _3691_/B _3691_/C vssd1 vssd1 vccd1 vccd1 _3707_/A sky130_fd_sc_hd__nand3_1
X_5430_ _5430_/A _5430_/B vssd1 vssd1 vccd1 vccd1 _5434_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5361_ _5351_/A _5351_/B _5349_/X vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__o21a_1
X_4312_ _4312_/A _4338_/A vssd1 vssd1 vccd1 vccd1 _4313_/B sky130_fd_sc_hd__or2_1
X_5292_ _5292_/A _5292_/B vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__and2_1
X_4243_ _4286_/A _4286_/B _4242_/X vssd1 vssd1 vccd1 vccd1 _4247_/B sky130_fd_sc_hd__a21o_2
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _5353_/A _4174_/B vssd1 vssd1 vccd1 vccd1 _4208_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3958_ _4989_/A _3958_/B vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3889_ _3889_/A _3889_/B vssd1 vssd1 vccd1 vccd1 _3890_/B sky130_fd_sc_hd__nand2_1
X_5628_ _5748_/A _5674_/A vssd1 vssd1 vccd1 vccd1 _5629_/A sky130_fd_sc_hd__nor2_1
X_5559_ _5679_/B _5559_/B vssd1 vssd1 vccd1 vccd1 _5564_/B sky130_fd_sc_hd__and2_1
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6396_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6518__100 vssd1 vssd1 vccd1 vccd1 _6518__100/HI _6626_/A sky130_fd_sc_hd__conb_1
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4930_ _4931_/A _4931_/B _4931_/C vssd1 vssd1 vccd1 vccd1 _4981_/S sky130_fd_sc_hd__o21ai_2
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4861_ _4861_/A _4861_/B _4861_/C vssd1 vssd1 vccd1 vccd1 _4866_/A sky130_fd_sc_hd__and3_1
X_6600_ _6600_/A _3295_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_3812_ _3812_/A _3846_/B vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__xnor2_1
X_4792_ _4918_/B _4792_/B vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3743_ _4905_/A _4904_/A vssd1 vssd1 vccd1 vccd1 _3743_/Y sky130_fd_sc_hd__nor2_1
X_3674_ _4830_/A _3718_/C vssd1 vssd1 vccd1 vccd1 _3703_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5413_ _5411_/Y _5413_/B vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__and2b_1
X_6393_ _6401_/CLK _6393_/D vssd1 vssd1 vccd1 vccd1 _6393_/Q sky130_fd_sc_hd__dfxtp_1
X_5344_ _5344_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _5348_/B sky130_fd_sc_hd__xnor2_2
XFILLER_114_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6467__49 vssd1 vssd1 vccd1 vccd1 _6467__49/HI _6572_/A sky130_fd_sc_hd__conb_1
X_5275_ _5275_/A _5275_/B vssd1 vssd1 vccd1 vccd1 _5275_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4226_ _4956_/A vssd1 vssd1 vccd1 vccd1 _4404_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4157_ _4177_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4157_/X sky130_fd_sc_hd__and2_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4088_ _4079_/C _4086_/Y _4089_/A _4087_/X vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__a211oi_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6481__63 vssd1 vssd1 vccd1 vccd1 _6481__63/HI _6589_/A sky130_fd_sc_hd__conb_1
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ _6331_/Q vssd1 vssd1 vccd1 vccd1 _3653_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5060_ _5060_/A _5353_/B vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__nand2_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4011_ _4213_/C vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5962_ _5962_/A vssd1 vssd1 vccd1 vccd1 _6323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4913_ _4867_/B _4913_/B vssd1 vssd1 vccd1 vccd1 _4913_/X sky130_fd_sc_hd__and2b_1
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5893_ _6424_/Q vssd1 vssd1 vccd1 vccd1 _5893_/Y sky130_fd_sc_hd__inv_2
X_4844_ _4847_/B _4847_/A vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4775_ _4775_/A _4798_/A vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__or2_1
X_3726_ _3726_/A _3726_/B vssd1 vssd1 vccd1 vccd1 _3735_/C sky130_fd_sc_hd__or2_1
X_3657_ _3657_/A _3657_/B vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__xnor2_2
X_3588_ _3588_/A _3588_/B vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__xnor2_1
X_6376_ _6396_/CLK _6376_/D vssd1 vssd1 vccd1 vccd1 _6376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5327_ _5327_/A _5327_/B vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5258_ _5258_/A _5266_/A vssd1 vssd1 vccd1 vccd1 _5259_/C sky130_fd_sc_hd__xnor2_1
X_4209_ _4246_/A _4246_/B vssd1 vssd1 vccd1 vccd1 _4209_/X sky130_fd_sc_hd__or2b_1
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5189_ _5100_/A _5196_/B _5184_/B _5183_/A vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__a31o_1
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4560_/A _4560_/B vssd1 vssd1 vccd1 vccd1 _4562_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3511_ _3511_/A _3511_/B vssd1 vssd1 vccd1 vccd1 _3519_/B sky130_fd_sc_hd__xor2_1
X_4491_ _4491_/A vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__inv_2
X_3442_ _3442_/A _3442_/B vssd1 vssd1 vccd1 vccd1 _3444_/B sky130_fd_sc_hd__nor2_1
X_6230_ _6393_/Q _6232_/B vssd1 vssd1 vccd1 vccd1 _6231_/A sky130_fd_sc_hd__and2_1
X_3373_ _5006_/A vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__clkbuf_2
X_6161_ _6161_/A vssd1 vssd1 vccd1 vccd1 _6367_/D sky130_fd_sc_hd__clkbuf_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5112_/A _5115_/B vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__xor2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6437__19 vssd1 vssd1 vccd1 vccd1 _6437__19/HI _6542_/A sky130_fd_sc_hd__conb_1
X_6092_ _6092_/A _6093_/A vssd1 vssd1 vccd1 vccd1 _6092_/X sky130_fd_sc_hd__or2b_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5044_/A _5040_/B _5041_/A _5039_/A vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__a31o_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5945_ _5945_/A _5950_/B vssd1 vssd1 vccd1 vccd1 _5946_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5876_ _5866_/X _5767_/X _5769_/Y _5823_/C vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4827_ _4813_/B _4807_/B _4807_/C vssd1 vssd1 vccd1 vccd1 _4832_/B sky130_fd_sc_hd__a21o_1
X_4758_ _4874_/A _4758_/B _4770_/A _4758_/D vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__and4_1
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4689_ _4682_/A _4769_/B _4687_/X _4723_/A vssd1 vssd1 vccd1 vccd1 _4706_/B sky130_fd_sc_hd__a22o_1
X_3709_ _3704_/A _3704_/B _3708_/X vssd1 vssd1 vccd1 vccd1 _3711_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6359_ _6361_/CLK _6359_/D vssd1 vssd1 vccd1 vccd1 _6359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6451__33 vssd1 vssd1 vccd1 vccd1 _6451__33/HI _6556_/A sky130_fd_sc_hd__conb_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _3991_/A _3978_/A vssd1 vssd1 vccd1 vccd1 _3992_/C sky130_fd_sc_hd__or2b_1
XFILLER_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5730_ _5730_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5730_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5661_ _5736_/B _5662_/B vssd1 vssd1 vccd1 vccd1 _5726_/B sky130_fd_sc_hd__nand2_1
X_5592_ _5592_/A _5592_/B vssd1 vssd1 vccd1 vccd1 _5593_/C sky130_fd_sc_hd__xor2_1
X_4612_ _4514_/A _4514_/B _4610_/X _4611_/X vssd1 vssd1 vccd1 vccd1 _5776_/B sky130_fd_sc_hd__a2bb2oi_1
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4543_ _5851_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4474_ _4474_/A _4474_/B _4474_/C vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__nand3_1
X_6213_ _6387_/Q _6213_/B vssd1 vssd1 vccd1 vccd1 _6214_/A sky130_fd_sc_hd__and2_1
X_3425_ _4651_/A _3406_/B _3395_/B _4711_/B vssd1 vssd1 vccd1 vccd1 _3426_/B sky130_fd_sc_hd__a22oi_1
X_6144_ _6144_/A vssd1 vssd1 vccd1 vccd1 _6361_/D sky130_fd_sc_hd__clkbuf_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3356_/A vssd1 vssd1 vccd1 vccd1 _3409_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3287_ _3291_/A vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__inv_2
X_6075_ _6083_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__and2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5083_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5928_ _5926_/A _5927_/Y _5928_/S vssd1 vssd1 vccd1 vccd1 _5929_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5859_ input8/X vssd1 vssd1 vccd1 vccd1 _6126_/B sky130_fd_sc_hd__inv_2
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4190_ _5316_/A _4135_/B _4424_/B _4189_/Y vssd1 vssd1 vccd1 vccd1 _4191_/C sky130_fd_sc_hd__a31oi_1
X_3210_ _3334_/A vssd1 vssd1 vccd1 vccd1 _3342_/A sky130_fd_sc_hd__buf_8
XFILLER_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _3974_/A vssd1 vssd1 vccd1 vccd1 _5095_/A sky130_fd_sc_hd__clkbuf_2
X_5713_ _4905_/C _5662_/B _5710_/Y _5916_/A _5829_/A vssd1 vssd1 vccd1 vccd1 _5714_/B
+ sky130_fd_sc_hd__o221a_1
X_5644_ _5681_/A _5803_/A vssd1 vssd1 vccd1 vccd1 _5644_/Y sky130_fd_sc_hd__xnor2_1
X_5575_ _5652_/A _5652_/B _5574_/X vssd1 vssd1 vccd1 vccd1 _5655_/B sky130_fd_sc_hd__a21o_1
XFILLER_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4526_ _5789_/A vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__inv_2
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4457_ _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__and2_1
X_3408_ _3424_/A _3441_/A vssd1 vssd1 vccd1 vccd1 _3421_/A sky130_fd_sc_hd__and2_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4388_ _4388_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__nor2_1
X_6127_ _6127_/A vssd1 vssd1 vccd1 vccd1 _6355_/D sky130_fd_sc_hd__clkbuf_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3339_/A vssd1 vssd1 vccd1 vccd1 _3339_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6058_ _6339_/Q _6036_/X _6057_/Y _6015_/X vssd1 vssd1 vccd1 vccd1 _6339_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5009_ _5009_/A _5009_/B _5009_/C vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__nor3_1
XFILLER_54_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _3690_/A _3706_/A _3690_/C vssd1 vssd1 vccd1 vccd1 _3691_/C sky130_fd_sc_hd__or3_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5360_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5379_/B sky130_fd_sc_hd__xor2_2
X_5291_ _5297_/C _5291_/B vssd1 vssd1 vccd1 vccd1 _5330_/B sky130_fd_sc_hd__xnor2_2
X_4311_ _4312_/A _4338_/A vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__nand2_1
X_4242_ _4241_/A _4242_/B vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4173_ _4173_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__xor2_1
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _3948_/A _3948_/B _3948_/C vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3888_ _4482_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _3888_/X sky130_fd_sc_hd__or2_1
X_5627_ _5627_/A _5627_/B vssd1 vssd1 vccd1 vccd1 _5674_/A sky130_fd_sc_hd__xnor2_4
X_5558_ _5693_/A _5692_/A _5557_/C vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__a21o_1
X_4509_ _4509_/A _4509_/B vssd1 vssd1 vccd1 vccd1 _4510_/B sky130_fd_sc_hd__nand2_2
X_5489_ _5545_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5498_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4839_/A _4838_/B _4838_/C vssd1 vssd1 vccd1 vccd1 _4861_/C sky130_fd_sc_hd__a21o_1
XFILLER_82_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3811_ _5684_/A _3858_/B _3822_/B _3810_/Y vssd1 vssd1 vccd1 vccd1 _3846_/B sky130_fd_sc_hd__a31o_1
XFILLER_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4791_ _4791_/A _4791_/B vssd1 vssd1 vccd1 vccd1 _4792_/B sky130_fd_sc_hd__xnor2_1
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3742_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3673_ _4755_/B vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__buf_2
X_5412_ _5413_/B _5411_/Y vssd1 vssd1 vccd1 vccd1 _5435_/B sky130_fd_sc_hd__or2b_1
X_6392_ _6396_/CLK _6392_/D vssd1 vssd1 vccd1 vccd1 _6392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _5338_/A _5337_/B _5337_/A vssd1 vssd1 vccd1 vccd1 _5348_/A sky130_fd_sc_hd__o21ba_2
XFILLER_114_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5274_ _5274_/A _5274_/B vssd1 vssd1 vccd1 vccd1 _5292_/A sky130_fd_sc_hd__nor2_1
X_4225_ _4225_/A _4225_/B vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__or2_2
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4087_ _4044_/X _4084_/X _4074_/Y _4082_/X vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4989_ _4989_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5061_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4010_ _4010_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _4213_/C sky130_fd_sc_hd__xor2_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5961_ _5959_/X _5961_/B vssd1 vssd1 vccd1 vccd1 _5962_/A sky130_fd_sc_hd__and2b_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _4951_/B _4951_/C _4951_/A vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__a21bo_2
X_5892_ _5743_/X _5891_/X _5870_/X _5851_/X vssd1 vssd1 vccd1 vccd1 _5892_/X sky130_fd_sc_hd__a2bb2o_1
X_4843_ _4404_/A _4820_/B _4837_/B _4842_/Y vssd1 vssd1 vccd1 vccd1 _4847_/A sky130_fd_sc_hd__a31o_2
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4774_ _4769_/Y _4772_/X _4775_/A _4773_/Y vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__a211oi_1
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3725_ _4891_/B _3494_/B _3718_/D _4891_/A vssd1 vssd1 vccd1 vccd1 _3726_/B sky130_fd_sc_hd__a22oi_1
X_3656_ _4828_/B _3656_/B vssd1 vssd1 vccd1 vccd1 _3681_/A sky130_fd_sc_hd__xnor2_2
X_3587_ _3587_/A _3587_/B vssd1 vssd1 vccd1 vccd1 _3637_/A sky130_fd_sc_hd__nand2_1
X_6375_ _6396_/CLK _6375_/D vssd1 vssd1 vccd1 vccd1 _6375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5326_ _5326_/A _5326_/B vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5257_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__nand2_1
X_4208_ _4208_/A _4208_/B vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__xor2_1
XFILLER_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _5188_/A _5188_/B vssd1 vssd1 vccd1 vccd1 _5192_/B sky130_fd_sc_hd__xor2_1
XFILLER_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4139_ _5322_/A _4169_/C vssd1 vssd1 vccd1 vccd1 _4140_/C sky130_fd_sc_hd__and2_1
XFILLER_95_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3510_ _3515_/A _3515_/B vssd1 vssd1 vccd1 vccd1 _3519_/A sky130_fd_sc_hd__xor2_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4490_ _4523_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__or2_1
XFILLER_109_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3441_ _3441_/A _3441_/B _3441_/C vssd1 vssd1 vccd1 vccd1 _3442_/B sky130_fd_sc_hd__and3_1
X_3372_ _5000_/A vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6160_ _6366_/Q _6164_/B vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__and2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5118_/A _5297_/B _5155_/B _5110_/Y vssd1 vssd1 vccd1 vccd1 _5115_/B sky130_fd_sc_hd__a31o_1
XFILLER_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6078_/A _6078_/C _6083_/C _6090_/X _6078_/B vssd1 vssd1 vccd1 vccd1 _6093_/A
+ sky130_fd_sc_hd__a311oi_4
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5087_/A _5087_/B _5087_/C vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__o21ai_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5944_/A vssd1 vssd1 vccd1 vccd1 _5950_/B sky130_fd_sc_hd__clkbuf_2
X_5875_ _5918_/A _5870_/A _5874_/X _5868_/A vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__o2bb2a_1
X_4826_ _4826_/A _4826_/B vssd1 vssd1 vccd1 vccd1 _4841_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4757_ _3646_/A _4855_/B _4855_/C _4895_/C _6332_/Q vssd1 vssd1 vccd1 vccd1 _4758_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4688_ _4780_/A _4688_/B _4872_/B _4728_/B vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__nand4_2
X_3708_ _3708_/A _3726_/A vssd1 vssd1 vccd1 vccd1 _3708_/X sky130_fd_sc_hd__or2_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3639_ _3617_/A _3617_/B _3625_/B vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__a21oi_2
X_6358_ _6361_/CLK _6358_/D vssd1 vssd1 vccd1 vccd1 _6358_/Q sky130_fd_sc_hd__dfxtp_1
X_5309_ _5625_/A _5625_/B _5625_/C vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6289_ _6416_/Q _6415_/Q _6289_/C vssd1 vssd1 vccd1 vccd1 _6290_/B sky130_fd_sc_hd__and3_1
XFILLER_102_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _5168_/A vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5660_ _5660_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__xor2_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4611_ _4611_/A _4611_/B vssd1 vssd1 vccd1 vccd1 _4611_/X sky130_fd_sc_hd__or2_1
X_5591_ _5591_/A _5591_/B vssd1 vssd1 vccd1 vccd1 _5593_/B sky130_fd_sc_hd__nor2_1
X_4542_ _4601_/B _4592_/B _4592_/C vssd1 vssd1 vccd1 vccd1 _4542_/X sky130_fd_sc_hd__a21o_1
X_4473_ _4495_/B _4496_/A _4496_/B _4472_/X vssd1 vssd1 vccd1 vccd1 _4594_/C sky130_fd_sc_hd__a31o_2
X_3424_ _3424_/A _3424_/B vssd1 vssd1 vccd1 vccd1 _3438_/A sky130_fd_sc_hd__and2_1
X_6212_ _6212_/A vssd1 vssd1 vccd1 vccd1 _6387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6143_ _6360_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6144_/A sky130_fd_sc_hd__and2_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _6346_/Q vssd1 vssd1 vccd1 vccd1 _3356_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3286_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3291_/A sky130_fd_sc_hd__buf_6
X_6074_ _6074_/A _6074_/B vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__or2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5025_ _5100_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5083_/B sky130_fd_sc_hd__nand2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5927_ _5927_/A _5927_/B vssd1 vssd1 vccd1 vccd1 _5927_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5858_ _6417_/Q _5858_/B vssd1 vssd1 vccd1 vccd1 _5858_/Y sky130_fd_sc_hd__nand2_1
X_4809_ _4809_/A _4760_/X vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__or2b_1
X_5789_ _5789_/A _5789_/B vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6511__93 vssd1 vssd1 vccd1 vccd1 _6511__93/HI _6619_/A sky130_fd_sc_hd__conb_1
XFILLER_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _5248_/A _3973_/B _3973_/C vssd1 vssd1 vccd1 vccd1 _3991_/A sky130_fd_sc_hd__and3_1
X_5712_ _5712_/A vssd1 vssd1 vccd1 vccd1 _5829_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5643_ _5730_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5643_/Y sky130_fd_sc_hd__nand2_1
X_5574_ _5484_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4525_ _4525_/A _4525_/B vssd1 vssd1 vccd1 vccd1 _4525_/X sky130_fd_sc_hd__or2_1
X_4456_ _4533_/A _4533_/B _4455_/Y vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__a21o_2
X_3407_ _3407_/A _3407_/B _3426_/A vssd1 vssd1 vccd1 vccd1 _3424_/A sky130_fd_sc_hd__or3b_1
X_4387_ _5486_/A _4387_/B _4387_/C vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__and3_1
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3338_ _3339_/A vssd1 vssd1 vccd1 vccd1 _3338_/Y sky130_fd_sc_hd__inv_2
X_6126_ _6401_/Q _6126_/B vssd1 vssd1 vccd1 vccd1 _6127_/A sky130_fd_sc_hd__and2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3269_ _3272_/A vssd1 vssd1 vccd1 vccd1 _3269_/Y sky130_fd_sc_hd__inv_2
X_6057_ _6099_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6057_/Y sky130_fd_sc_hd__nand2_1
X_5008_ _5008_/A _5013_/C vssd1 vssd1 vccd1 vccd1 _5009_/C sky130_fd_sc_hd__xnor2_1
XFILLER_39_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5290_ _5290_/A _5290_/B vssd1 vssd1 vccd1 vccd1 _5291_/B sky130_fd_sc_hd__nand2_1
X_4310_ _5371_/A _5441_/C _4336_/A vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__and3_1
X_4241_ _4241_/A _4242_/B vssd1 vssd1 vccd1 vccd1 _4286_/B sky130_fd_sc_hd__xnor2_1
X_4172_ _5290_/A _4221_/B vssd1 vssd1 vccd1 vccd1 _4173_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3956_ _4493_/A _3956_/B vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__nor2_2
XFILLER_23_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5626_ _5626_/A _5626_/B vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__nor2_2
X_3887_ _3887_/A _3887_/B _3887_/C vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__and3_1
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5557_ _5693_/A _5692_/A _5557_/C vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__nand3_1
X_4508_ _4159_/Y _4167_/A _4127_/B _4129_/X vssd1 vssd1 vccd1 vccd1 _4509_/B sky130_fd_sc_hd__a211o_1
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5488_ _5488_/A _5511_/A vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__xnor2_1
X_4439_ _4445_/A _4445_/B _4446_/B vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__or3_1
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _4782_/A _4782_/B _4789_/Y vssd1 vssd1 vccd1 vccd1 _4918_/B sky130_fd_sc_hd__a21bo_1
X_3810_ _3810_/A _3810_/B vssd1 vssd1 vccd1 vccd1 _3810_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3741_ _3741_/A _3741_/B vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__or2_2
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3672_ _3672_/A _3699_/A _3699_/C _3699_/D vssd1 vssd1 vccd1 vccd1 _3683_/B sky130_fd_sc_hd__nand4_2
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5411_ _5411_/A _5411_/B vssd1 vssd1 vccd1 vccd1 _5411_/Y sky130_fd_sc_hd__xnor2_1
X_6391_ _6396_/CLK _6391_/D vssd1 vssd1 vccd1 vccd1 _6391_/Q sky130_fd_sc_hd__dfxtp_1
X_5342_ _5344_/A _5344_/B vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__or2b_1
XFILLER_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5273_ _5198_/A _5240_/B _5240_/C vssd1 vssd1 vccd1 vccd1 _5274_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ _4109_/A _4412_/B _4191_/C vssd1 vssd1 vccd1 vccd1 _4225_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4155_ _4161_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__xor2_1
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4086_ _4122_/B vssd1 vssd1 vccd1 vccd1 _4086_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4988_ _5169_/B vssd1 vssd1 vccd1 vccd1 _5335_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3939_ _4140_/B vssd1 vssd1 vccd1 vccd1 _4317_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5609_ _5609_/A _5609_/B vssd1 vssd1 vccd1 vccd1 _5615_/A sky130_fd_sc_hd__nand2_2
X_6589_ _6589_/A _3281_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6472__54 vssd1 vssd1 vccd1 vccd1 _6472__54/HI _6577_/A sky130_fd_sc_hd__conb_1
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5960_ _5933_/B _5956_/X _5957_/Y _3354_/X vssd1 vssd1 vccd1 vccd1 _5961_/B sky130_fd_sc_hd__a31o_1
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _3364_/B _5748_/X _5750_/X _5871_/X vssd1 vssd1 vccd1 vccd1 _5891_/X sky130_fd_sc_hd__o22a_1
X_4911_ _4882_/A _4909_/A _4866_/B _4868_/X vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__a211o_1
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _4842_/A _4842_/B vssd1 vssd1 vccd1 vccd1 _4842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _4768_/A _4768_/C _4768_/B vssd1 vssd1 vccd1 vccd1 _4773_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _4895_/B vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__clkbuf_2
X_3655_ _3655_/A _3655_/B vssd1 vssd1 vccd1 vccd1 _3669_/A sky130_fd_sc_hd__xor2_2
X_3586_ _3586_/A _3586_/B vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__nand2_1
X_6374_ _6388_/CLK _6374_/D vssd1 vssd1 vccd1 vccd1 _6374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5325_ _5325_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__xor2_2
X_5256_ _5168_/A _5101_/B _5250_/B _5249_/B vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__a31o_1
X_4207_ _4207_/A _4207_/B vssd1 vssd1 vccd1 vccd1 _4465_/B sky130_fd_sc_hd__xnor2_2
X_5187_ _5188_/B _5188_/A vssd1 vssd1 vccd1 vccd1 _5191_/B sky130_fd_sc_hd__or2b_1
XFILLER_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4138_ _4095_/A _4140_/B _4347_/B _5281_/A vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__a22oi_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4069_ _4069_/A _4069_/B _5287_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__or4bb_1
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3440_ _3440_/A _3440_/B _3447_/A vssd1 vssd1 vccd1 vccd1 _3482_/A sky130_fd_sc_hd__or3_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3371_ _4989_/A vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__buf_2
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5110_ _5110_/A _5160_/A vssd1 vssd1 vccd1 vccd1 _5110_/Y sky130_fd_sc_hd__nor2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6343_/Q _6074_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5041_/B vssd1 vssd1 vccd1 vccd1 _5087_/C sky130_fd_sc_hd__xnor2_1
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5943_ _5940_/A _5940_/B _5938_/A vssd1 vssd1 vccd1 vccd1 _5946_/A sky130_fd_sc_hd__o21ai_2
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5874_ _5866_/A _5775_/Y _5779_/Y _5871_/X vssd1 vssd1 vccd1 vccd1 _5874_/X sky130_fd_sc_hd__o2bb2a_1
X_4825_ _4825_/A _4825_/B vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__xnor2_2
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4756_ _4756_/A _4855_/B _4855_/C _4874_/C vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__nand4_1
X_4687_ _4780_/A _4872_/B _4728_/B _4688_/B vssd1 vssd1 vccd1 vccd1 _4687_/X sky130_fd_sc_hd__a22o_1
X_3707_ _3707_/A _3707_/B _3730_/A vssd1 vssd1 vccd1 vccd1 _3712_/A sky130_fd_sc_hd__nand3_2
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3638_ _3640_/B _3640_/A vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__or2b_1
X_6426_ _6426_/CLK _6426_/D vssd1 vssd1 vccd1 vccd1 _6426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6357_ _6361_/CLK _6357_/D vssd1 vssd1 vccd1 vccd1 _6357_/Q sky130_fd_sc_hd__dfxtp_1
X_3569_ _4659_/B vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5308_ _5310_/A _5310_/B vssd1 vssd1 vccd1 vccd1 _5625_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6288_ _6415_/Q _6289_/C _6287_/Y vssd1 vssd1 vccd1 vccd1 _6415_/D sky130_fd_sc_hd__o21a_1
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5239_ _5244_/B _5239_/B vssd1 vssd1 vccd1 vccd1 _5240_/C sky130_fd_sc_hd__and2b_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6442__24 vssd1 vssd1 vccd1 vccd1 _6442__24/HI _6547_/A sky130_fd_sc_hd__conb_1
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4610_ _4611_/A _4611_/B _4525_/X _4609_/X vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__a22o_1
X_5590_ _5148_/B _5590_/B vssd1 vssd1 vccd1 vccd1 _5593_/A sky130_fd_sc_hd__and2b_1
X_4541_ _5950_/A _4543_/B _4540_/X vssd1 vssd1 vccd1 vccd1 _4592_/C sky130_fd_sc_hd__o21ai_1
X_4472_ _4472_/A _4472_/B _4472_/C vssd1 vssd1 vccd1 vccd1 _4472_/X sky130_fd_sc_hd__and3_1
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3423_ _3407_/A _3407_/B _3426_/A vssd1 vssd1 vccd1 vccd1 _3424_/B sky130_fd_sc_hd__o21bai_1
X_6211_ _6386_/Q _6213_/B vssd1 vssd1 vccd1 vccd1 _6212_/A sky130_fd_sc_hd__and2_1
X_6142_ _6142_/A vssd1 vssd1 vccd1 vccd1 _6360_/D sky130_fd_sc_hd__clkbuf_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _5672_/A vssd1 vssd1 vccd1 vccd1 _3354_/X sky130_fd_sc_hd__buf_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3285_ input1/X vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__clkbuf_4
X_6073_ _6074_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6083_/A sky130_fd_sc_hd__nand2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5024_ _5096_/B vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5926_ _5926_/A _5944_/A vssd1 vssd1 vccd1 vccd1 _5927_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5857_ _5847_/Y _5852_/X _5853_/Y _5856_/Y vssd1 vssd1 vccd1 vccd1 _5857_/X sky130_fd_sc_hd__a211o_1
X_4808_ _4808_/A _4832_/A vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__nand2_1
X_5788_ _5796_/B _5788_/B vssd1 vssd1 vccd1 vccd1 _5788_/Y sky130_fd_sc_hd__nor2_1
X_4739_ _4739_/A _4739_/B _4739_/C vssd1 vssd1 vccd1 vccd1 _4740_/B sky130_fd_sc_hd__and3_1
XFILLER_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6409_ _6425_/CLK _6409_/D vssd1 vssd1 vccd1 vccd1 _6409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _5288_/A vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _5711_/A vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5642_ _5796_/A _5688_/A vssd1 vssd1 vccd1 vccd1 _5730_/B sky130_fd_sc_hd__xor2_1
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5573_ _5660_/A _5660_/B _5572_/X vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__a21o_2
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4524_ _4520_/Y _4522_/Y _4523_/X vssd1 vssd1 vccd1 vccd1 _4525_/B sky130_fd_sc_hd__a21boi_1
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4455_ _4455_/A _4455_/B vssd1 vssd1 vccd1 vccd1 _4455_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3406_ _4711_/B _3406_/B _3406_/C vssd1 vssd1 vccd1 vccd1 _3426_/A sky130_fd_sc_hd__and3_1
X_4386_ _4388_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _4387_/C sky130_fd_sc_hd__nor2_1
XFILLER_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3337_ _3339_/A vssd1 vssd1 vccd1 vccd1 _3337_/Y sky130_fd_sc_hd__inv_2
X_6125_ _6125_/A vssd1 vssd1 vccd1 vccd1 _6354_/D sky130_fd_sc_hd__clkbuf_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3268_ _3272_/A vssd1 vssd1 vccd1 vccd1 _3268_/Y sky130_fd_sc_hd__inv_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6056_/A _6056_/B vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5007_ _5007_/A _5007_/B vssd1 vssd1 vccd1 vccd1 _5013_/C sky130_fd_sc_hd__xor2_2
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5909_ _5954_/A vssd1 vssd1 vccd1 vccd1 _5909_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4240_ _4238_/A _4238_/B _4239_/X vssd1 vssd1 vccd1 vccd1 _4242_/B sky130_fd_sc_hd__o21ai_2
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4171_ _5287_/A _4302_/B _4180_/A _4169_/X vssd1 vssd1 vccd1 vccd1 _4173_/A sky130_fd_sc_hd__a31o_2
XFILLER_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3955_ _3954_/B _3955_/B vssd1 vssd1 vccd1 vccd1 _3956_/B sky130_fd_sc_hd__and2b_1
X_5625_ _5625_/A _5625_/B _5625_/C vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__and3_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3886_ _3854_/A _3854_/B _3848_/B _3848_/A vssd1 vssd1 vccd1 vccd1 _3887_/C sky130_fd_sc_hd__a211o_1
X_5556_ _5556_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _5557_/C sky130_fd_sc_hd__xor2_1
X_4507_ _4515_/A _4515_/B _4468_/X vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__a21oi_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5487_ _5487_/A _5487_/B vssd1 vssd1 vccd1 vccd1 _5511_/A sky130_fd_sc_hd__nand2_2
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _4441_/A _4441_/C _4441_/B vssd1 vssd1 vccd1 vccd1 _4446_/B sky130_fd_sc_hd__a21boi_1
X_6478__60 vssd1 vssd1 vccd1 vccd1 _6478__60/HI _6586_/A sky130_fd_sc_hd__conb_1
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4369_ _4369_/A _4369_/B vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__or2_1
XFILLER_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6134_/A input5/X vssd1 vssd1 vccd1 vccd1 _6109_/A sky130_fd_sc_hd__and2_1
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6039_ _6040_/A _6040_/B vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__and2_1
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6525__107 vssd1 vssd1 vccd1 vccd1 _6525__107/HI _6633_/A sky130_fd_sc_hd__conb_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3740_ _4814_/A _3589_/A _3718_/D _4891_/B vssd1 vssd1 vccd1 vccd1 _3741_/B sky130_fd_sc_hd__a22oi_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3671_ _6330_/Q _3671_/B vssd1 vssd1 vccd1 vccd1 _4851_/A sky130_fd_sc_hd__and2_2
X_5410_ _5373_/B _5406_/Y _5440_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5413_/B sky130_fd_sc_hd__o22ai_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6390_ _6396_/CLK _6390_/D vssd1 vssd1 vccd1 vccd1 _6390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5341_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5344_/B sky130_fd_sc_hd__xor2_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5272_ _5272_/A _5272_/B vssd1 vssd1 vccd1 vccd1 _5307_/B sky130_fd_sc_hd__xnor2_2
X_4223_ _4223_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__xnor2_1
X_4154_ _5335_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__nand2_1
X_4085_ _4074_/Y _4082_/X _4044_/X _4084_/X vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__a211oi_2
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _4987_/A _4987_/B vssd1 vssd1 vccd1 vccd1 _5169_/B sky130_fd_sc_hd__xnor2_2
X_3938_ _3938_/A _3938_/B vssd1 vssd1 vccd1 vccd1 _4140_/B sky130_fd_sc_hd__xor2_4
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3869_ _3808_/A _3875_/A _3817_/Y vssd1 vssd1 vccd1 vccd1 _3870_/B sky130_fd_sc_hd__o21ba_1
XFILLER_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6588_ _6588_/A _3280_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
X_5608_ _5608_/A _5608_/B vssd1 vssd1 vccd1 vccd1 _5609_/B sky130_fd_sc_hd__or2_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5539_ _5539_/A _5539_/B vssd1 vssd1 vccd1 vccd1 _5544_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _5883_/X _5886_/X _5889_/X vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__a21o_1
X_4910_ _4953_/B _4953_/C _4953_/A vssd1 vssd1 vccd1 vccd1 _4951_/C sky130_fd_sc_hd__a21bo_1
X_4841_ _4841_/A _4841_/B vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__xor2_4
X_4772_ _4785_/C _4772_/B vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__xor2_1
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3723_ _4904_/A _3729_/A _3723_/C vssd1 vssd1 vccd1 vccd1 _3735_/B sky130_fd_sc_hd__nand3_1
X_3654_ _3651_/A _3652_/A _3651_/B _3656_/B _4828_/B vssd1 vssd1 vccd1 vccd1 _3670_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3585_ _3585_/A _3585_/B vssd1 vssd1 vccd1 vccd1 _3600_/B sky130_fd_sc_hd__xor2_2
X_6373_ _6388_/CLK _6373_/D vssd1 vssd1 vccd1 vccd1 _6373_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6388_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5324_ _5324_/A _5392_/B vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5255_ _5255_/A vssd1 vssd1 vccd1 vccd1 _5350_/B sky130_fd_sc_hd__clkbuf_4
X_4206_ _4206_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _4207_/B sky130_fd_sc_hd__xor2_1
X_6448__30 vssd1 vssd1 vccd1 vccd1 _6448__30/HI _6553_/A sky130_fd_sc_hd__conb_1
X_5186_ _5219_/B _5219_/C _5219_/A vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__a21bo_1
XFILLER_110_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4135_/A _4135_/B _4182_/A vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__a21oi_2
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4068_ _4095_/A _4068_/B _4068_/C vssd1 vssd1 vccd1 vccd1 _4069_/B sky130_fd_sc_hd__and3_2
XFILLER_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3370_ _5102_/A vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__buf_2
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5100_/A _5040_/B vssd1 vssd1 vccd1 vccd1 _5041_/B sky130_fd_sc_hd__nand2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5942_ _5936_/A _5909_/X _5941_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _6320_/D sky130_fd_sc_hd__o211a_1
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5873_ _5785_/X _5870_/X _5872_/X _4634_/X vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__o2bb2a_1
X_4824_ _4824_/A _4824_/B _4824_/C vssd1 vssd1 vccd1 vccd1 _4967_/B sky130_fd_sc_hd__nand3_2
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4755_ _4762_/A _4755_/B _4755_/C vssd1 vssd1 vccd1 vccd1 _4874_/C sky130_fd_sc_hd__and3b_1
X_3706_ _3706_/A _3706_/B _3706_/C vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__nand3_2
X_4686_ _4802_/B vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__clkbuf_2
X_3637_ _3637_/A _3637_/B vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__xor2_1
X_6425_ _6425_/CLK _6425_/D vssd1 vssd1 vccd1 vccd1 _6425_/Q sky130_fd_sc_hd__dfxtp_1
X_3568_ _3653_/A vssd1 vssd1 vccd1 vccd1 _3612_/A sky130_fd_sc_hd__clkbuf_2
X_6356_ _6401_/CLK _6356_/D vssd1 vssd1 vccd1 vccd1 _6356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5307_ _5307_/A _5307_/B vssd1 vssd1 vccd1 vccd1 _5310_/B sky130_fd_sc_hd__xnor2_2
X_3499_ _3570_/C vssd1 vssd1 vccd1 vccd1 _3718_/D sky130_fd_sc_hd__clkbuf_2
X_6287_ _6304_/A _6287_/B vssd1 vssd1 vccd1 vccd1 _6287_/Y sky130_fd_sc_hd__nor2_1
X_5238_ _4109_/A _5255_/A _5237_/Y vssd1 vssd1 vccd1 vccd1 _5239_/B sky130_fd_sc_hd__a21bo_1
X_5169_ _5248_/B _5169_/B vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__nand2_2
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4540_ _4540_/A _4540_/B vssd1 vssd1 vccd1 vccd1 _4540_/X sky130_fd_sc_hd__or2_1
X_4471_ _4165_/Y _4469_/Y _4470_/X vssd1 vssd1 vccd1 vccd1 _4496_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3422_ _3441_/B _3422_/B vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__and2_1
X_6210_ _6210_/A vssd1 vssd1 vccd1 vccd1 _6386_/D sky130_fd_sc_hd__clkbuf_1
X_6141_ _6359_/Q _6145_/B vssd1 vssd1 vccd1 vccd1 _6142_/A sky130_fd_sc_hd__and2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _5044_/A vssd1 vssd1 vccd1 vccd1 _5672_/A sky130_fd_sc_hd__clkbuf_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3284_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__inv_2
X_6072_ _6074_/B vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__clkbuf_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5087_/A _5023_/B vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__or2_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5925_ _5937_/B vssd1 vssd1 vccd1 vccd1 _5944_/A sky130_fd_sc_hd__clkbuf_2
X_5856_ _6417_/Q _5858_/B vssd1 vssd1 vccd1 vccd1 _5856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4807_ _4813_/B _4807_/B _4807_/C vssd1 vssd1 vccd1 vccd1 _4832_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5787_ _5787_/A _5787_/B vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__nor2_1
X_4738_ _4739_/A _4739_/B _4739_/C vssd1 vssd1 vccd1 vccd1 _4740_/A sky130_fd_sc_hd__a21oi_1
X_4669_ _4855_/B _4855_/C vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__and2_1
XFILLER_107_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408_ _6425_/CLK _6408_/D vssd1 vssd1 vccd1 vccd1 _6408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6339_ _6345_/CLK _6339_/D vssd1 vssd1 vccd1 vccd1 _6339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6502__84 vssd1 vssd1 vccd1 vccd1 _6502__84/HI _6610_/A sky130_fd_sc_hd__conb_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3971_ _5096_/A _3969_/X _3973_/C vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__a21oi_1
X_5710_ _5714_/A _5710_/B vssd1 vssd1 vccd1 vccd1 _5710_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5641_ _5738_/A _5695_/A vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__and2b_1
X_5572_ _5508_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5572_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4523_ _4523_/A _4523_/B _4554_/A vssd1 vssd1 vccd1 vccd1 _4523_/X sky130_fd_sc_hd__or3_1
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _4538_/A _4545_/A _4453_/X vssd1 vssd1 vccd1 vccd1 _4533_/B sky130_fd_sc_hd__o21ai_4
X_3405_ _4697_/B vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4385_ _5538_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _4386_/B sky130_fd_sc_hd__nor2_1
X_3336_ _3339_/A vssd1 vssd1 vccd1 vccd1 _3336_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6124_ _6353_/Q _6314_/B vssd1 vssd1 vccd1 vccd1 _6125_/A sky130_fd_sc_hd__and2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6049_/A _6049_/B _6047_/A vssd1 vssd1 vccd1 vccd1 _6056_/B sky130_fd_sc_hd__o21ai_1
X_5006_ _5006_/A _5168_/B vssd1 vssd1 vccd1 vccd1 _5007_/B sky130_fd_sc_hd__nand2_1
X_3267_ _3279_/A vssd1 vssd1 vccd1 vccd1 _3272_/A sky130_fd_sc_hd__buf_6
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5908_ _5933_/B vssd1 vssd1 vccd1 vccd1 _5954_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5839_ _3364_/A _5798_/X _5820_/X _5796_/Y vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4170_ _4140_/C _4168_/X _4169_/X vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__o21ba_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ _3955_/B _3954_/B vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__and2b_2
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3885_ _3925_/A _3925_/B vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__nor2_1
X_5624_ _5630_/A _5630_/B _5583_/Y vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5555_ _5547_/B _5554_/Y _5555_/C _5555_/D vssd1 vssd1 vccd1 vccd1 _5692_/A sky130_fd_sc_hd__and4bb_2
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5486_ _5486_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4506_ _5777_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _4506_/Y sky130_fd_sc_hd__nor2_1
X_4437_ _4573_/A _4440_/C _4188_/X vssd1 vssd1 vccd1 vccd1 _4441_/B sky130_fd_sc_hd__or3b_1
X_4368_ _4368_/A _4368_/B vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__xor2_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6294_/B _6107_/B vssd1 vssd1 vccd1 vccd1 _6346_/D sky130_fd_sc_hd__nor2_1
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4299_ _4314_/A _4314_/B _4298_/X vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__a21o_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3319_/Y sky130_fd_sc_hd__inv_2
X_6493__75 vssd1 vssd1 vccd1 vccd1 _6493__75/HI _6601_/A sky130_fd_sc_hd__conb_1
X_6038_ _6038_/A _6046_/B vssd1 vssd1 vccd1 vccd1 _6040_/B sky130_fd_sc_hd__xor2_1
XFILLER_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3670_ _3670_/A _3670_/B vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__xor2_4
X_5340_ _5358_/A _5358_/B _5339_/X vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__o21ba_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5271_ _5271_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5625_/A sky130_fd_sc_hd__xnor2_2
X_4222_ _4244_/A _4244_/B vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__xor2_1
X_4153_ _4160_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__xnor2_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _4047_/B _4044_/C _4083_/Y _4027_/X vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4986_ _5067_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3937_ _3937_/A _3937_/B vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__xnor2_1
XFILLER_11_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ _3881_/A _3881_/B vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__xor2_1
X_3799_ _3843_/A _3799_/B vssd1 vssd1 vccd1 vccd1 _3800_/C sky130_fd_sc_hd__nor2_1
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5607_ _5608_/A _5608_/B vssd1 vssd1 vccd1 vccd1 _5609_/A sky130_fd_sc_hd__nand2_1
X_6587_ _6587_/A _3278_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5538_ _5538_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5539_/B sky130_fd_sc_hd__or2_1
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5469_ _5471_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__nand2_1
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4840_ _4841_/B _4841_/A vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__and2b_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4771_ _4905_/A _4812_/B vssd1 vssd1 vccd1 vccd1 _4772_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3722_ _3722_/A vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__buf_2
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3653_ _3653_/A _3671_/B vssd1 vssd1 vccd1 vccd1 _4828_/B sky130_fd_sc_hd__nand2_4
X_6372_ _6388_/CLK _6372_/D vssd1 vssd1 vccd1 vccd1 _6372_/Q sky130_fd_sc_hd__dfxtp_1
X_5323_ _5333_/A _5351_/A vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__xor2_2
X_3584_ _3577_/A _3577_/B _3587_/B vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__a21bo_2
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5254_ _5262_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _5272_/A sky130_fd_sc_hd__xnor2_2
X_4205_ _4468_/B _4205_/B vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__xnor2_4
X_5185_ _5175_/A _5175_/B _5174_/Y vssd1 vssd1 vccd1 vccd1 _5219_/A sky130_fd_sc_hd__o21bai_1
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4136_ _5406_/A _4213_/D _4136_/C vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__and3_1
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6463__45 vssd1 vssd1 vccd1 vccd1 _6463__45/HI _6568_/A sky130_fd_sc_hd__conb_1
X_4067_ _4095_/A _4068_/B _4068_/C vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__a21oi_2
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ _5055_/A _5055_/B _5092_/A _5092_/B vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__or4_2
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6639_ _6639_/A _3332_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5941_ _5954_/A _5941_/B vssd1 vssd1 vccd1 vccd1 _5941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5872_ _5866_/X _5788_/Y _5790_/Y _5871_/X vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__o2bb2a_1
X_4823_ _4825_/A _4825_/B vssd1 vssd1 vccd1 vccd1 _4824_/C sky130_fd_sc_hd__nand2_1
X_4754_ _4776_/A _4754_/B _4754_/C vssd1 vssd1 vccd1 vccd1 _4768_/A sky130_fd_sc_hd__or3_1
X_3705_ _3705_/A _3705_/B _3705_/C vssd1 vssd1 vccd1 vccd1 _3706_/C sky130_fd_sc_hd__nand3_1
X_4685_ _4777_/A _4777_/B _4684_/X vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__a21oi_1
X_3636_ _3655_/A _3655_/B _3635_/X vssd1 vssd1 vccd1 vccd1 _3640_/B sky130_fd_sc_hd__o21a_1
X_6508__90 vssd1 vssd1 vccd1 vccd1 _6508__90/HI _6616_/A sky130_fd_sc_hd__conb_1
X_6424_ _6425_/CLK _6424_/D vssd1 vssd1 vccd1 vccd1 _6424_/Q sky130_fd_sc_hd__dfxtp_1
X_3567_ _4659_/B _3646_/C _3570_/C _3653_/A vssd1 vssd1 vccd1 vccd1 _3573_/A sky130_fd_sc_hd__a22o_1
X_6355_ _6401_/CLK _6355_/D vssd1 vssd1 vccd1 vccd1 _6355_/Q sky130_fd_sc_hd__dfxtp_1
X_5306_ _5136_/A _5317_/B _5301_/B _5305_/X vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__a31o_2
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6286_ _6415_/Q _6289_/C vssd1 vssd1 vccd1 vccd1 _6287_/B sky130_fd_sc_hd__and2_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5237_ _5237_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5237_/Y sky130_fd_sc_hd__nand2_1
X_3498_ _3607_/A vssd1 vssd1 vccd1 vccd1 _3570_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5168_ _5168_/A _5168_/B vssd1 vssd1 vccd1 vccd1 _5172_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4119_ _5257_/A _4118_/B _4118_/C _4118_/D vssd1 vssd1 vccd1 vccd1 _4121_/C sky130_fd_sc_hd__a22o_1
X_5099_ _5711_/A _5214_/B _5114_/B _5098_/Y vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__a31o_1
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _4470_/A _4470_/B _4470_/C vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__or3_2
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3421_ _3421_/A _3421_/B vssd1 vssd1 vccd1 vccd1 _3422_/B sky130_fd_sc_hd__or2_1
X_3352_ _5100_/A vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6140_ _6140_/A vssd1 vssd1 vccd1 vccd1 _6359_/D sky130_fd_sc_hd__clkbuf_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3283_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6071_ _6341_/Q _6036_/X _6070_/X _5948_/X vssd1 vssd1 vccd1 vccd1 _6341_/D sky130_fd_sc_hd__o211a_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5021_/B _5022_/B vssd1 vssd1 vccd1 vccd1 _5023_/B sky130_fd_sc_hd__and2b_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6433__15 vssd1 vssd1 vccd1 vccd1 _6433__15/HI _6538_/A sky130_fd_sc_hd__conb_1
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _5829_/A _5917_/B _5915_/X vssd1 vssd1 vccd1 vccd1 _5927_/A sky130_fd_sc_hd__a21o_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5855_ _3354_/X _5825_/X _5854_/X _5743_/X vssd1 vssd1 vccd1 vccd1 _5858_/B sky130_fd_sc_hd__o2bb2a_1
X_4806_ _4808_/A _4806_/B _4806_/C vssd1 vssd1 vccd1 vccd1 _4807_/C sky130_fd_sc_hd__and3_1
X_5786_ _5766_/B _5775_/A _5758_/A _5766_/A vssd1 vssd1 vccd1 vccd1 _5787_/B sky130_fd_sc_hd__o211a_1
X_4737_ _4934_/A _4934_/B vssd1 vssd1 vccd1 vccd1 _4739_/C sky130_fd_sc_hd__xnor2_1
X_4668_ _4668_/A _4747_/A vssd1 vssd1 vccd1 vccd1 _4684_/B sky130_fd_sc_hd__nand2_1
X_3619_ _4895_/B vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__clkbuf_2
X_6407_ _6425_/CLK _6407_/D vssd1 vssd1 vccd1 vccd1 _6407_/Q sky130_fd_sc_hd__dfxtp_1
X_4599_ _4604_/A _4604_/B _4598_/X vssd1 vssd1 vccd1 vccd1 _4599_/X sky130_fd_sc_hd__a21bo_1
XFILLER_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6338_ _6345_/CLK _6338_/D vssd1 vssd1 vccd1 vccd1 _6338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6269_ _6280_/A _6269_/B vssd1 vssd1 vccd1 vccd1 _6269_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6499__81 vssd1 vssd1 vccd1 vccd1 _6499__81/HI _6607_/A sky130_fd_sc_hd__conb_1
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _5198_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _3973_/C sky130_fd_sc_hd__and2_1
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5640_ _5640_/A _5640_/B vssd1 vssd1 vccd1 vccd1 _5695_/A sky130_fd_sc_hd__xor2_4
XFILLER_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5571_ _5529_/Y _5664_/B _5663_/A vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__a21o_2
X_4522_ _4523_/A _4523_/B _4554_/A vssd1 vssd1 vccd1 vccd1 _4522_/Y sky130_fd_sc_hd__o21ai_1
X_4453_ _4453_/A _4421_/A vssd1 vssd1 vccd1 vccd1 _4453_/X sky130_fd_sc_hd__or2b_1
XFILLER_104_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3404_ _4673_/B vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ _5691_/A _4573_/B vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6123_ _6123_/A vssd1 vssd1 vccd1 vccd1 _6353_/D sky130_fd_sc_hd__clkbuf_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _3339_/A vssd1 vssd1 vccd1 vccd1 _3335_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3266_ _3266_/A vssd1 vssd1 vccd1 vccd1 _3266_/Y sky130_fd_sc_hd__inv_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6052_/X _6054_/B vssd1 vssd1 vccd1 vccd1 _6056_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5005_ _5064_/A _5113_/B vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__nand2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5907_ _5928_/S vssd1 vssd1 vccd1 vccd1 _5933_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5838_ _6412_/Q _5824_/Y _5827_/X _6413_/Q _5837_/X vssd1 vssd1 vccd1 vccd1 _5838_/X
+ sky130_fd_sc_hd__a221o_1
X_5769_ _5769_/A _5769_/B vssd1 vssd1 vccd1 vccd1 _5769_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _3953_/A _3953_/B vssd1 vssd1 vccd1 vccd1 _3954_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3884_ _3882_/A _3882_/B _3890_/A vssd1 vssd1 vccd1 vccd1 _3925_/B sky130_fd_sc_hd__o21a_1
X_5623_ _5736_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _5766_/B sky130_fd_sc_hd__and2_1
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5554_ _5362_/A _5560_/B _4441_/A vssd1 vssd1 vccd1 vccd1 _5554_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5485_ _5485_/A _5485_/B vssd1 vssd1 vccd1 vccd1 _5508_/A sky130_fd_sc_hd__xnor2_2
X_4505_ _4618_/A _4512_/B vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__or2_1
X_4436_ _6316_/Q _4436_/B vssd1 vssd1 vccd1 vccd1 _4440_/C sky130_fd_sc_hd__nand2_1
X_4367_ _5441_/C vssd1 vssd1 vccd1 vccd1 _5471_/C sky130_fd_sc_hd__clkbuf_2
X_3318_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3318_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6106_/A _6106_/B vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__xor2_1
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4298_ _5387_/A _4298_/B _4298_/C vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__and3_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _6027_/X _6029_/X _6030_/X _6028_/Y vssd1 vssd1 vccd1 vccd1 _6046_/B sky130_fd_sc_hd__o22a_2
X_3249_ _3253_/A vssd1 vssd1 vccd1 vccd1 _3249_/Y sky130_fd_sc_hd__inv_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6469__51 vssd1 vssd1 vccd1 vccd1 _6469__51/HI _6574_/A sky130_fd_sc_hd__conb_1
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _5225_/B _5229_/X _5265_/Y _5269_/Y vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__o211ai_2
X_4221_ _5392_/A _4221_/B vssd1 vssd1 vccd1 vccd1 _4244_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _5297_/A _4152_/B vssd1 vssd1 vccd1 vccd1 _4160_/B sky130_fd_sc_hd__nand2_1
X_4083_ _4027_/A _4027_/B _4027_/C vssd1 vssd1 vccd1 vccd1 _4083_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _5121_/B vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3936_ _5000_/A _4174_/B vssd1 vssd1 vccd1 vccd1 _3937_/A sky130_fd_sc_hd__nand2_1
X_3867_ _5067_/A _4041_/B vssd1 vssd1 vccd1 vccd1 _3881_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3798_ _3810_/B _3798_/B vssd1 vssd1 vccd1 vccd1 _3799_/B sky130_fd_sc_hd__and2_1
X_6586_ _6586_/A _3277_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
X_5606_ _5606_/A _5606_/B vssd1 vssd1 vccd1 vccd1 _5608_/B sky130_fd_sc_hd__and2_1
XFILLER_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5537_ _5537_/A _5537_/B vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__or2_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5468_ _5468_/A _5468_/B vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__xor2_2
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4419_ _4419_/A _4419_/B vssd1 vssd1 vccd1 vccd1 _4451_/B sky130_fd_sc_hd__nor2_1
X_5399_ _5399_/A _5399_/B vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__xor2_2
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6531__113 vssd1 vssd1 vccd1 vccd1 _6531__113/HI _6639_/A sky130_fd_sc_hd__conb_1
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4770_ _4770_/A _4770_/B vssd1 vssd1 vccd1 vccd1 _4785_/C sky130_fd_sc_hd__nand2_1
X_3721_ _3729_/A _3723_/C _3722_/A vssd1 vssd1 vccd1 vccd1 _3735_/A sky130_fd_sc_hd__a21o_1
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3652_ _3652_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3656_/B sky130_fd_sc_hd__xnor2_2
X_3583_ _3586_/A _3586_/B vssd1 vssd1 vccd1 vccd1 _3587_/B sky130_fd_sc_hd__or2_1
X_6371_ _6388_/CLK _6371_/D vssd1 vssd1 vccd1 vccd1 _6371_/Q sky130_fd_sc_hd__dfxtp_1
X_5322_ _5322_/A _5322_/B vssd1 vssd1 vccd1 vccd1 _5351_/A sky130_fd_sc_hd__nand2_2
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5253_ _5253_/A _5253_/B vssd1 vssd1 vccd1 vccd1 _5262_/B sky130_fd_sc_hd__or2_1
X_4204_ _4207_/A _4202_/X _4203_/X vssd1 vssd1 vccd1 vccd1 _4205_/B sky130_fd_sc_hd__o21a_2
X_5184_ _5184_/A _5184_/B vssd1 vssd1 vccd1 vccd1 _5219_/C sky130_fd_sc_hd__xnor2_1
X_4135_ _4135_/A _4135_/B vssd1 vssd1 vccd1 vccd1 _4136_/C sky130_fd_sc_hd__xor2_1
XFILLER_110_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4066_ _5317_/A _4066_/B vssd1 vssd1 vccd1 vccd1 _4068_/C sky130_fd_sc_hd__and2_1
XFILLER_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _4968_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _5092_/B sky130_fd_sc_hd__xnor2_4
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3919_ _3917_/A _3917_/B _3951_/A vssd1 vssd1 vccd1 vccd1 _3921_/B sky130_fd_sc_hd__a21o_1
X_4899_ _4899_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6638_ _6638_/A _3333_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_6569_ _6569_/A _3257_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6439__21 vssd1 vssd1 vccd1 vccd1 _6439__21/HI _6544_/A sky130_fd_sc_hd__conb_1
XFILLER_105_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5940_ _5940_/A _5940_/B vssd1 vssd1 vccd1 vccd1 _5941_/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5871_ _5871_/A _5871_/B _5817_/A vssd1 vssd1 vccd1 vccd1 _5871_/X sky130_fd_sc_hd__or3b_2
X_4822_ _4822_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4825_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4753_ _4779_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4754_/C sky130_fd_sc_hd__xnor2_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3704_ _3704_/A _3704_/B vssd1 vssd1 vccd1 vccd1 _3706_/B sky130_fd_sc_hd__xnor2_1
X_4684_ _4680_/B _4684_/B vssd1 vssd1 vccd1 vccd1 _4684_/X sky130_fd_sc_hd__and2b_1
X_6423_ _6423_/CLK _6423_/D vssd1 vssd1 vccd1 vccd1 _6423_/Q sky130_fd_sc_hd__dfxtp_1
X_3635_ _3635_/A _3634_/B vssd1 vssd1 vccd1 vccd1 _3635_/X sky130_fd_sc_hd__or2b_1
X_6354_ _6401_/CLK _6354_/D vssd1 vssd1 vccd1 vccd1 _6354_/Q sky130_fd_sc_hd__dfxtp_1
X_3566_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3646_/C sky130_fd_sc_hd__clkbuf_2
X_5305_ _5300_/A _5305_/B vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__and2b_1
X_6285_ _6414_/Q _6280_/B _6284_/Y vssd1 vssd1 vccd1 vccd1 _6414_/D sky130_fd_sc_hd__o21a_1
X_3497_ _3356_/A _3359_/A _6338_/Q vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__a21o_1
X_5236_ _5236_/A vssd1 vssd1 vccd1 vccd1 _5317_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5175_/A _5167_/B vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4118_ _5257_/A _4118_/B _4118_/C _4118_/D vssd1 vssd1 vccd1 vccd1 _4121_/B sky130_fd_sc_hd__nand4_4
X_5098_ _5137_/A _5178_/A vssd1 vssd1 vccd1 vccd1 _5098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4049_ _4050_/A _4049_/B _4049_/C vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__nand3_1
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3420_ _3441_/A _3441_/B _3441_/C vssd1 vssd1 vccd1 vccd1 _3442_/A sky130_fd_sc_hd__a21oi_1
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3351_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5100_/A sky130_fd_sc_hd__buf_2
XFILLER_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3282_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6070_ _6077_/B _6068_/Y _6069_/Y vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__a21o_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5021_ _5022_/B _5021_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__and2b_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5923_ _6100_/A vssd1 vssd1 vccd1 vccd1 _6134_/A sky130_fd_sc_hd__buf_2
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ _5818_/X _4619_/X _5849_/X _5742_/B vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__o2bb2a_1
X_4805_ _4805_/A _4805_/B _4805_/C _4830_/D vssd1 vssd1 vccd1 vccd1 _4806_/C sky130_fd_sc_hd__or4b_1
X_5785_ _5785_/A vssd1 vssd1 vccd1 vccd1 _5785_/X sky130_fd_sc_hd__clkbuf_2
X_4736_ _4931_/B _4736_/B vssd1 vssd1 vccd1 vccd1 _4934_/B sky130_fd_sc_hd__or2_1
X_4667_ _4763_/A _4873_/B _4668_/A _4667_/D vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__nand4_1
X_6406_ _6425_/CLK _6406_/D vssd1 vssd1 vccd1 vccd1 _6406_/Q sky130_fd_sc_hd__dfxtp_1
X_3618_ _6326_/Q vssd1 vssd1 vccd1 vccd1 _4895_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4598_ _5777_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4598_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6337_ _6345_/CLK _6337_/D vssd1 vssd1 vccd1 vccd1 _6337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3549_ _3588_/A _3588_/B vssd1 vssd1 vccd1 vccd1 _3553_/C sky130_fd_sc_hd__nand2_1
X_6268_ _6408_/Q _6407_/Q _6268_/C vssd1 vssd1 vccd1 vccd1 _6269_/B sky130_fd_sc_hd__and3_1
X_5219_ _5219_/A _5219_/B _5219_/C vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__and3_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6199_ _6380_/Q _6379_/Q _6382_/Q _6381_/Q vssd1 vssd1 vccd1 vccd1 _6199_/X sky130_fd_sc_hd__and4_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5570_ _5570_/A _5570_/B vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__nor2_1
X_4521_ _4521_/A _4521_/B vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__xnor2_4
X_4452_ _4544_/B _4553_/A _4544_/A vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__o21ai_4
X_3403_ _4659_/B vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__clkbuf_2
X_4383_ _4383_/A _5532_/B _4383_/C vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__and3_1
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6122_ _6352_/Q _6314_/B vssd1 vssd1 vccd1 vccd1 _6123_/A sky130_fd_sc_hd__and2_1
X_3334_ _3334_/A vssd1 vssd1 vccd1 vccd1 _3339_/A sky130_fd_sc_hd__buf_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3265_ _3266_/A vssd1 vssd1 vccd1 vccd1 _3265_/Y sky130_fd_sc_hd__inv_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6339_/Q _6059_/A vssd1 vssd1 vccd1 vccd1 _6054_/B sky130_fd_sc_hd__or2_1
X_5004_ _5004_/A _5004_/B vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__nand2_2
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5906_ _5902_/X _5903_/Y _5904_/X _5905_/X vssd1 vssd1 vccd1 vccd1 _5928_/S sky130_fd_sc_hd__o22a_1
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5837_ _6412_/Q _5824_/Y _5834_/X _5836_/X vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__o22a_1
X_5768_ _4506_/Y _5776_/A _5776_/B _5778_/A vssd1 vssd1 vccd1 vccd1 _5769_/B sky130_fd_sc_hd__o31a_1
XFILLER_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4719_ _4722_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4723_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5699_ _5699_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5700_/A sky130_fd_sc_hd__or2_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3952_ _3997_/B _3997_/C _3997_/A vssd1 vssd1 vccd1 vccd1 _3955_/B sky130_fd_sc_hd__a21boi_1
X_3883_ _3889_/A _3889_/B vssd1 vssd1 vccd1 vccd1 _3890_/A sky130_fd_sc_hd__or2_1
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5622_ _5622_/A _5622_/B vssd1 vssd1 vccd1 vccd1 _5736_/B sky130_fd_sc_hd__xor2_4
X_5553_ _5553_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _5693_/A sky130_fd_sc_hd__xnor2_2
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4504_ _4535_/A _4535_/B vssd1 vssd1 vccd1 vccd1 _4512_/B sky130_fd_sc_hd__and2_1
X_5484_ _5484_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__xnor2_4
XFILLER_117_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4435_ _5518_/A vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__inv_2
XFILLER_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _4366_/A _4366_/B vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__xor2_4
X_3317_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3317_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6103_/X _6104_/X _6041_/A vssd1 vssd1 vccd1 vccd1 _6106_/B sky130_fd_sc_hd__a21bo_1
X_4297_ _4297_/A _4298_/C vssd1 vssd1 vccd1 vccd1 _4314_/B sky130_fd_sc_hd__xnor2_2
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3248_/A vssd1 vssd1 vccd1 vccd1 _3253_/A sky130_fd_sc_hd__buf_12
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6484__66 vssd1 vssd1 vccd1 vccd1 _6484__66/HI _6592_/A sky130_fd_sc_hd__conb_1
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4220_ _5428_/A vssd1 vssd1 vccd1 vccd1 _5392_/A sky130_fd_sc_hd__buf_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4151_ _4141_/A _4143_/B _4141_/B vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__o21ba_1
X_4082_ _4122_/A _4122_/B _4122_/C _4122_/D vssd1 vssd1 vccd1 vccd1 _4082_/X sky130_fd_sc_hd__or4_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4984_ _5180_/B vssd1 vssd1 vccd1 vccd1 _5121_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _3920_/B _3918_/B _3918_/C vssd1 vssd1 vccd1 vccd1 _3951_/B sky130_fd_sc_hd__a21oi_1
XFILLER_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3866_ _5122_/A vssd1 vssd1 vccd1 vccd1 _5067_/A sky130_fd_sc_hd__buf_2
X_5605_ _5605_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5608_/A sky130_fd_sc_hd__xnor2_1
X_6585_ _6585_/A _3276_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_3797_ _5028_/A _3858_/B vssd1 vssd1 vccd1 vccd1 _3798_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5536_ _5492_/A _5535_/B _5535_/C vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5467_ _5467_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__xnor2_1
X_4418_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4419_/B sky130_fd_sc_hd__and2_1
X_5398_ _5398_/A _5398_/B vssd1 vssd1 vccd1 vccd1 _5419_/B sky130_fd_sc_hd__xor2_2
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4349_ _4349_/A _4349_/B vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__xnor2_1
XFILLER_86_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6019_ _4630_/A _6001_/S _6017_/X _6018_/Y _6282_/A vssd1 vssd1 vccd1 vccd1 _6019_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3720_ _3720_/A _3720_/B _3741_/A vssd1 vssd1 vccd1 vccd1 _3723_/C sky130_fd_sc_hd__nand3_1
X_3651_ _3651_/A _3651_/B vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__nand2_1
X_3582_ _4745_/A _3716_/D _3650_/B _4855_/A vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__a22o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6370_ _6388_/CLK _6370_/D vssd1 vssd1 vccd1 vccd1 _6370_/Q sky130_fd_sc_hd__dfxtp_1
X_5321_ _5350_/A _5428_/B vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5252_ _5252_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _5253_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4203_ _4206_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _4203_/X sky130_fd_sc_hd__or2_1
X_5183_ _5183_/A _5183_/B vssd1 vssd1 vccd1 vccd1 _5184_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4134_ _5367_/A vssd1 vssd1 vccd1 vccd1 _5406_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4212_/A vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4967_ _4915_/Y _4967_/B vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__and2b_1
XFILLER_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3918_ _3920_/B _3918_/B _3918_/C vssd1 vssd1 vccd1 vccd1 _3951_/A sky130_fd_sc_hd__and3_1
X_4898_ _4904_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _4902_/C sky130_fd_sc_hd__nor2_1
X_3849_ _5044_/A _3849_/B vssd1 vssd1 vccd1 vccd1 _3849_/Y sky130_fd_sc_hd__nand2_1
X_6637_ _6637_/A _3335_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_6568_ _6568_/A _3256_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5519_ _5519_/A _5519_/B vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__xnor2_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6454__36 vssd1 vssd1 vccd1 vccd1 _6454__36/HI _6559_/A sky130_fd_sc_hd__conb_1
XFILLER_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5870_/A vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4821_ _5967_/A _4924_/B _4816_/B _4820_/X vssd1 vssd1 vccd1 vccd1 _4825_/A sky130_fd_sc_hd__a31o_1
X_4752_ _4752_/A _4780_/C vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__xor2_1
X_4683_ _4683_/A _4683_/B vssd1 vssd1 vccd1 vccd1 _4777_/B sky130_fd_sc_hd__xnor2_1
X_3703_ _3722_/A _3703_/B vssd1 vssd1 vccd1 vccd1 _3704_/B sky130_fd_sc_hd__nor2_1
X_3634_ _3635_/A _3634_/B vssd1 vssd1 vccd1 vccd1 _3655_/B sky130_fd_sc_hd__xor2_2
X_6422_ _6423_/CLK _6422_/D vssd1 vssd1 vccd1 vccd1 _6422_/Q sky130_fd_sc_hd__dfxtp_1
X_3565_ _3565_/A _3565_/B vssd1 vssd1 vccd1 vccd1 _3603_/A sky130_fd_sc_hd__xnor2_1
X_6353_ _6401_/CLK _6353_/D vssd1 vssd1 vccd1 vccd1 _6353_/Q sky130_fd_sc_hd__dfxtp_1
X_3496_ _4765_/D _3494_/X _3507_/A vssd1 vssd1 vccd1 vccd1 _3506_/A sky130_fd_sc_hd__a21bo_1
X_5304_ _5307_/B _5307_/A vssd1 vssd1 vccd1 vccd1 _5625_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6284_ _6304_/A _6289_/C vssd1 vssd1 vccd1 vccd1 _6284_/Y sky130_fd_sc_hd__nor2_1
X_5235_ _5455_/B _5455_/C vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__and2_1
XFILLER_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5166_ _5166_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5167_/B sky130_fd_sc_hd__nor2_1
X_4117_ _5297_/A _3969_/X _4096_/B _4114_/X vssd1 vssd1 vccd1 vccd1 _4118_/D sky130_fd_sc_hd__a211o_1
XFILLER_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5097_ _5137_/A _5178_/A vssd1 vssd1 vccd1 vccd1 _5114_/B sky130_fd_sc_hd__xor2_2
X_4048_ _3996_/X _4045_/Y _4027_/X _4044_/X vssd1 vssd1 vccd1 vccd1 _4049_/C sky130_fd_sc_hd__a211o_1
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _4627_/A _5997_/B _5998_/X vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__o21ai_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ _5211_/A vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__buf_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3281_/Y sky130_fd_sc_hd__inv_2
X_5020_ _5027_/B _5020_/B vssd1 vssd1 vccd1 vccd1 _5021_/B sky130_fd_sc_hd__xnor2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ _5765_/X _5909_/X _5919_/Y _5921_/X vssd1 vssd1 vccd1 vccd1 _6317_/D sky130_fd_sc_hd__o211a_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5853_ _6415_/Q _5844_/Y _5852_/X _5847_/Y vssd1 vssd1 vccd1 vccd1 _5853_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4804_ _3612_/A _4895_/C _4850_/B _3647_/A vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__a22o_1
X_5784_ _5784_/A _5784_/B _5784_/C _5783_/Y vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__or4b_1
X_4735_ _4924_/A _4820_/B _4734_/C vssd1 vssd1 vccd1 vccd1 _4736_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4666_ _3647_/A _4694_/A _4663_/A _4895_/C _4745_/A vssd1 vssd1 vccd1 vccd1 _4667_/D
+ sky130_fd_sc_hd__a32o_1
X_3617_ _3617_/A _3617_/B vssd1 vssd1 vccd1 vccd1 _3624_/A sky130_fd_sc_hd__xnor2_1
X_4597_ _4614_/A _4614_/B _4596_/C vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__o21ai_1
X_6405_ _6425_/CLK _6405_/D vssd1 vssd1 vccd1 vccd1 _6405_/Q sky130_fd_sc_hd__dfxtp_1
X_3548_ _3548_/A _3548_/B vssd1 vssd1 vccd1 vccd1 _3588_/B sky130_fd_sc_hd__xnor2_1
X_6336_ _6345_/CLK _6336_/D vssd1 vssd1 vccd1 vccd1 _6336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3479_ _3479_/A _3479_/B vssd1 vssd1 vccd1 vccd1 _3480_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6267_ _6407_/Q _6268_/C _6266_/Y vssd1 vssd1 vccd1 vccd1 _6407_/D sky130_fd_sc_hd__o21a_1
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5218_ _5219_/A _5219_/B _5219_/C vssd1 vssd1 vccd1 vccd1 _5218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6198_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6382_/D sky130_fd_sc_hd__clkbuf_1
X_5149_ _5591_/A _5591_/B vssd1 vssd1 vccd1 vccd1 _5596_/A sky130_fd_sc_hd__xnor2_4
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4520_ _5790_/A _4562_/A vssd1 vssd1 vccd1 vccd1 _4520_/Y sky130_fd_sc_hd__nor2_1
X_4451_ _4451_/A _4451_/B vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__xor2_2
X_3402_ _6330_/Q vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4382_ _4404_/A _6319_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _5532_/B sky130_fd_sc_hd__and3_2
X_6121_ _6121_/A vssd1 vssd1 vccd1 vccd1 _6352_/D sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3333_/A vssd1 vssd1 vccd1 vccd1 _3333_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3264_ _3266_/A vssd1 vssd1 vccd1 vccd1 _3264_/Y sky130_fd_sc_hd__inv_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6339_/Q _6059_/A vssd1 vssd1 vccd1 vccd1 _6052_/X sky130_fd_sc_hd__and2_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5003_ _4995_/A _4995_/B _4979_/C _4979_/D vssd1 vssd1 vccd1 vccd1 _5004_/B sky130_fd_sc_hd__o22ai_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5905_ _6356_/Q _6365_/Q vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__and2b_1
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5836_ _6273_/A _5831_/X _5828_/X vssd1 vssd1 vccd1 vccd1 _5836_/X sky130_fd_sc_hd__o21a_1
X_5767_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5767_/X sky130_fd_sc_hd__and2_1
XFILLER_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4718_ _4724_/A _4724_/B vssd1 vssd1 vccd1 vccd1 _4722_/B sky130_fd_sc_hd__xnor2_1
X_5698_ _5706_/A _5698_/B vssd1 vssd1 vccd1 vccd1 _5699_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4649_ _4745_/B vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6319_ _6361_/CLK _6319_/D vssd1 vssd1 vccd1 vccd1 _6319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _3951_/A _3951_/B _3949_/X vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__or3b_1
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3882_ _3882_/A _3882_/B vssd1 vssd1 vccd1 vccd1 _3889_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5621_ _5634_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5736_/A sky130_fd_sc_hd__and2b_1
X_5552_ _5556_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__nand2_1
X_4503_ _4165_/Y _4469_/Y _4496_/A _4470_/X vssd1 vssd1 vccd1 vccd1 _4535_/B sky130_fd_sc_hd__o211ai_4
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _5485_/A _5485_/B _5482_/X vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__a21o_2
X_4434_ _5546_/A _4188_/X _4436_/B _5514_/A vssd1 vssd1 vccd1 vccd1 _4441_/C sky130_fd_sc_hd__a22o_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4365_ _5392_/A _4109_/B _4374_/B _4364_/X vssd1 vssd1 vccd1 vccd1 _4380_/A sky130_fd_sc_hd__a31o_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _3334_/A vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__buf_12
X_6104_ _6104_/A _6104_/B _6103_/B _6093_/A vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__or4bb_1
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4296_ _5471_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4298_/C sky130_fd_sc_hd__and2_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6040_/A _6032_/X _6034_/Y vssd1 vssd1 vccd1 vccd1 _6336_/D sky130_fd_sc_hd__a21oi_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3247_/A vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5819_ _6106_/A _6104_/A _5848_/A vssd1 vssd1 vccd1 vccd1 _5868_/C sky130_fd_sc_hd__nor3_1
XFILLER_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4150_ _4156_/B _4156_/A vssd1 vssd1 vccd1 vccd1 _4150_/X sky130_fd_sc_hd__and2b_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4081_ _4075_/A _4075_/B _4075_/C vssd1 vssd1 vccd1 vccd1 _4122_/D sky130_fd_sc_hd__a21oi_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _4979_/C _5004_/A _4983_/C _4983_/D vssd1 vssd1 vccd1 vccd1 _5180_/B sky130_fd_sc_hd__and4b_2
XFILLER_17_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3934_ _3934_/A _3948_/A vssd1 vssd1 vccd1 vccd1 _3997_/B sky130_fd_sc_hd__or2b_1
X_3865_ _5096_/A vssd1 vssd1 vccd1 vccd1 _5122_/A sky130_fd_sc_hd__buf_2
XFILLER_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5604_ _4274_/A _5045_/B _5603_/X vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__o21ai_1
X_6584_ _6584_/A _3275_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
X_3796_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5535_ _5546_/A _5535_/B _5535_/C vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__and3_1
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5466_ _5466_/A _5466_/B vssd1 vssd1 vccd1 vccd1 _5494_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4417_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5397_ _5399_/A _5399_/B _5394_/A vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__o21ai_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _5297_/A _4109_/B _4341_/A _4347_/X vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__a31o_1
X_4279_ _4278_/B _4279_/B vssd1 vssd1 vccd1 vccd1 _4280_/B sky130_fd_sc_hd__and2b_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6018_ _5756_/A _6011_/X _5992_/X vssd1 vssd1 vccd1 vccd1 _6018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3650_ _3685_/A _3650_/B _4800_/C vssd1 vssd1 vccd1 vccd1 _3651_/B sky130_fd_sc_hd__nand3_1
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3581_ _6327_/Q vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__clkbuf_2
X_5320_ _5318_/A _5318_/B _5365_/A vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__o21ai_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _5294_/A _5294_/B _5245_/A vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__a21oi_2
X_4202_ _4206_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _4202_/X sky130_fd_sc_hd__and2_1
X_5182_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5183_/B sky130_fd_sc_hd__nor3_1
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4133_ _4272_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__and2_1
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4064_ _5102_/A _4347_/B _4100_/B _4062_/X vssd1 vssd1 vccd1 vccd1 _4071_/B sky130_fd_sc_hd__a31o_1
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4966_ _4950_/A _4950_/B _4916_/X vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3917_ _3917_/A _3917_/B vssd1 vssd1 vccd1 vccd1 _3918_/C sky130_fd_sc_hd__xor2_1
X_4897_ _4902_/B _4897_/B vssd1 vssd1 vccd1 vccd1 _4904_/B sky130_fd_sc_hd__or2_1
X_6636_ _6636_/A _3336_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_3848_ _3848_/A _3848_/B vssd1 vssd1 vccd1 vccd1 _3887_/B sky130_fd_sc_hd__nand2_1
X_6567_ _6567_/A _3253_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_3779_ _6322_/Q vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__clkbuf_2
X_5518_ _5518_/A _5546_/B vssd1 vssd1 vccd1 vccd1 _5519_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5449_ _5465_/A _5447_/Y _5448_/Y vssd1 vssd1 vccd1 vccd1 _5451_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4820_ _5979_/A _4820_/B _4820_/C vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__and3_1
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4672_/X _4755_/B _4751_/C vssd1 vssd1 vccd1 vccd1 _4780_/C sky130_fd_sc_hd__and3b_1
X_4682_ _4682_/A _4728_/B vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__nand2_1
X_3702_ _4874_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _3722_/A sky130_fd_sc_hd__nand2_1
X_6421_ _6423_/CLK _6421_/D vssd1 vssd1 vccd1 vccd1 _6421_/Q sky130_fd_sc_hd__dfxtp_1
X_3633_ _3657_/A _3657_/B _3631_/Y vssd1 vssd1 vccd1 vccd1 _3634_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3564_ _3564_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _3813_/A sky130_fd_sc_hd__nor2_2
X_6352_ _6401_/CLK _6352_/D vssd1 vssd1 vccd1 vccd1 _6352_/Q sky130_fd_sc_hd__dfxtp_1
X_5303_ _5295_/A _5295_/B _5302_/X vssd1 vssd1 vccd1 vccd1 _5307_/A sky130_fd_sc_hd__o21ai_2
X_3495_ _4756_/A _3494_/B _3466_/B _4765_/D vssd1 vssd1 vccd1 vccd1 _3507_/A sky130_fd_sc_hd__a22o_1
X_6283_ _6414_/Q _6413_/Q _6283_/C vssd1 vssd1 vccd1 vccd1 _6289_/C sky130_fd_sc_hd__and3_1
XFILLER_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _5234_/A _5492_/C vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__and2_1
X_5165_ _5166_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__and2_1
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _5290_/A vssd1 vssd1 vccd1 vccd1 _5297_/A sky130_fd_sc_hd__buf_2
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5096_ _5096_/A _5096_/B vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__nand2_2
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4047_ _4047_/A _4047_/B vssd1 vssd1 vccd1 vccd1 _4049_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6521__103 vssd1 vssd1 vccd1 vccd1 _6521__103/HI _6629_/A sky130_fd_sc_hd__conb_1
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5987_/A _5987_/B _5756_/C _5997_/B vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__a2bb2o_1
X_4949_ _4967_/B _4948_/C _4948_/A vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6619_ _6619_/A _3315_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
XFILLER_106_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6514__96 vssd1 vssd1 vccd1 vccd1 _6514__96/HI _6622_/A sky130_fd_sc_hd__conb_1
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3280_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3280_/Y sky130_fd_sc_hd__inv_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5921_ _6115_/B vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5852_ _5743_/X _5850_/X _5825_/X _5851_/X vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__a2bb2o_1
X_4803_ _4888_/A _4802_/B _4813_/A _4802_/D vssd1 vssd1 vccd1 vccd1 _4807_/B sky130_fd_sc_hd__a22o_1
X_5783_ _5783_/A _5783_/B vssd1 vssd1 vccd1 vccd1 _5783_/Y sky130_fd_sc_hd__nand2_1
X_4734_ _4924_/A _4820_/B _4734_/C vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__and3_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4665_ _6038_/A _3671_/B _4762_/A vssd1 vssd1 vccd1 vccd1 _4895_/C sky130_fd_sc_hd__o21ba_2
X_3616_ _4891_/A _3615_/X _3586_/B vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__a21boi_2
X_4596_ _4614_/A _4614_/B _4596_/C vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__or3_1
X_6404_ _6425_/CLK _6404_/D vssd1 vssd1 vccd1 vccd1 _6404_/Q sky130_fd_sc_hd__dfxtp_1
X_3547_ _3547_/A _3547_/B vssd1 vssd1 vccd1 vccd1 _3548_/A sky130_fd_sc_hd__nand2_1
X_6335_ _6396_/CLK _6335_/D vssd1 vssd1 vccd1 vccd1 _6335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3478_ _3479_/A _3479_/B vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6266_ _6280_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6266_/Y sky130_fd_sc_hd__nor2_1
X_5217_ _5264_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__or2b_1
XFILLER_69_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6197_ _6381_/Q _6213_/B vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__and2_1
XFILLER_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5148_ _5590_/B _5148_/B vssd1 vssd1 vccd1 vccd1 _5591_/B sky130_fd_sc_hd__xor2_4
X_5079_ _5079_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__nand2_1
XFILLER_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4450_ _4552_/B _4560_/A _4552_/A vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__a21oi_2
X_3401_ _3395_/A _3406_/B _3395_/B _4710_/A vssd1 vssd1 vccd1 vccd1 _3407_/B sky130_fd_sc_hd__a22oi_1
X_4381_ _4381_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__xnor2_4
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6120_ _6351_/Q _6314_/B vssd1 vssd1 vccd1 vccd1 _6121_/A sky130_fd_sc_hd__and2_1
X_3332_ _3333_/A vssd1 vssd1 vccd1 vccd1 _3332_/Y sky130_fd_sc_hd__inv_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3266_/A vssd1 vssd1 vccd1 vccd1 _3263_/Y sky130_fd_sc_hd__inv_2
X_6051_ _6338_/Q _6036_/X _6050_/Y _6015_/X vssd1 vssd1 vccd1 vccd1 _6338_/D sky130_fd_sc_hd__o211a_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5002_ _5064_/A _5040_/B _5065_/B vssd1 vssd1 vccd1 vccd1 _5009_/B sky130_fd_sc_hd__and3_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5904_ _6365_/Q _6356_/Q vssd1 vssd1 vccd1 vccd1 _5904_/X sky130_fd_sc_hd__and2b_1
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5835_ _6410_/Q vssd1 vssd1 vccd1 vccd1 _6273_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5766_ _5766_/A _5766_/B _5775_/A vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__or3_1
X_4717_ _4780_/A _4854_/B _4716_/X _4627_/A vssd1 vssd1 vccd1 vccd1 _4724_/B sky130_fd_sc_hd__a22oi_4
X_5697_ _5697_/A vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__buf_2
XFILLER_108_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648_ _4660_/B _4648_/B vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__xor2_2
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4579_ _4579_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__xnor2_4
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6318_ _6361_/CLK _6318_/D vssd1 vssd1 vccd1 vccd1 _6318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6249_ _6247_/X _6248_/X _6355_/D vssd1 vssd1 vccd1 vccd1 _6249_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ _3951_/A _3951_/B _3949_/X vssd1 vssd1 vccd1 vccd1 _3997_/C sky130_fd_sc_hd__o21bai_1
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ _3881_/A _3881_/B vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__or2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ _5666_/A _5666_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__and2_1
X_5551_ _5555_/C _5514_/B _5547_/B _5550_/X vssd1 vssd1 vccd1 vccd1 _5556_/B sky130_fd_sc_hd__a31o_1
X_4502_ _4496_/A _4470_/X _4165_/Y _4469_/Y vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__a211o_2
X_5482_ _5481_/B _5482_/B vssd1 vssd1 vccd1 vccd1 _5482_/X sky130_fd_sc_hd__and2b_1
X_4433_ _4433_/A _4433_/B vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__and2_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4364_ _4363_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4364_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4295_ _5424_/A _4391_/B _4391_/C vssd1 vssd1 vccd1 vccd1 _4314_/A sky130_fd_sc_hd__and3_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__inv_2
X_6103_ _6103_/A _6103_/B _6103_/C vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__or3_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3247_/A vssd1 vssd1 vccd1 vccd1 _3246_/Y sky130_fd_sc_hd__inv_2
X_6034_ _6040_/A _6036_/A _5911_/X vssd1 vssd1 vccd1 vccd1 _6034_/Y sky130_fd_sc_hd__o21ai_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5818_ _6106_/A _6104_/A _5848_/A vssd1 vssd1 vccd1 vccd1 _5818_/X sky130_fd_sc_hd__and3b_1
X_5749_ _5805_/A _5805_/B vssd1 vssd1 vccd1 vccd1 _5750_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4080_ _5214_/A _3858_/B _4079_/C _4079_/D vssd1 vssd1 vccd1 vccd1 _4122_/C sky130_fd_sc_hd__a22oi_4
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6475__57 vssd1 vssd1 vccd1 vccd1 _6475__57/HI _6583_/A sky130_fd_sc_hd__conb_1
XFILLER_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _4630_/A _4716_/X _4981_/X vssd1 vssd1 vccd1 vccd1 _4983_/D sky130_fd_sc_hd__a21oi_1
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3933_ _3933_/A _3934_/A _5068_/A _3903_/B vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__or4bb_1
X_3864_ _5288_/A vssd1 vssd1 vccd1 vccd1 _5096_/A sky130_fd_sc_hd__clkbuf_2
X_5603_ _5044_/A _5029_/B _5031_/A _5045_/A vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__a22o_1
X_3795_ _5211_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3810_/B sky130_fd_sc_hd__nand2_1
X_6583_ _6583_/A _3274_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
X_5534_ _5424_/A _5471_/B _5532_/B _5549_/A vssd1 vssd1 vccd1 vccd1 _5535_/C sky130_fd_sc_hd__a31o_1
XFILLER_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5465_ _5465_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__xnor2_2
X_4416_ _4422_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4418_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5396_ _5433_/A _5555_/D vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__nand2_1
X_4347_ _5392_/A _4347_/B _4347_/C vssd1 vssd1 vccd1 vccd1 _4347_/X sky130_fd_sc_hd__and3_1
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4278_ _4279_/B _4278_/B vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__and2b_1
X_3229_ _3229_/A vssd1 vssd1 vccd1 vccd1 _3229_/Y sky130_fd_sc_hd__inv_2
X_6017_ _5756_/A _4629_/A _6004_/X _6010_/B vssd1 vssd1 vccd1 vccd1 _6017_/X sky130_fd_sc_hd__a31o_1
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _3671_/B vssd1 vssd1 vccd1 vccd1 _3716_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5250_ _5250_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__xnor2_2
X_4201_ _4197_/X _4201_/B vssd1 vssd1 vccd1 vccd1 _4206_/B sky130_fd_sc_hd__and2b_1
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5181_ _5182_/A _5182_/B _5182_/C vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__o21a_1
XFILLER_96_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _4231_/A vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4016_/B _4061_/Y _4062_/X vssd1 vssd1 vccd1 vccd1 _4100_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _5106_/A _5106_/B vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__nand2_2
XFILLER_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3916_ _3915_/A _3915_/B _3992_/B _5697_/A vssd1 vssd1 vccd1 vccd1 _3918_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4896_ _4895_/A _4956_/B _4891_/D _3685_/A vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__a22oi_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6635_ _6635_/A _3337_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_3847_ _3847_/A vssd1 vssd1 vccd1 vccd1 _3848_/B sky130_fd_sc_hd__inv_2
X_3778_ _4041_/B vssd1 vssd1 vccd1 vccd1 _3849_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6566_ _6566_/A _3252_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
X_5517_ _5517_/A _5517_/B vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5448_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5448_/Y sky130_fd_sc_hd__nor2_1
X_5379_ _5378_/B _5379_/B vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6445__27 vssd1 vssd1 vccd1 vccd1 _6445__27/HI _6550_/A sky130_fd_sc_hd__conb_1
XFILLER_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _4756_/A _4850_/B vssd1 vssd1 vccd1 vccd1 _4752_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4681_ _4711_/D vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__clkbuf_2
X_3701_ _4805_/B vssd1 vssd1 vccd1 vccd1 _4886_/B sky130_fd_sc_hd__clkbuf_2
X_6420_ _6425_/CLK _6420_/D vssd1 vssd1 vccd1 vccd1 _6420_/Q sky130_fd_sc_hd__dfxtp_1
X_3632_ _3593_/B _3660_/A _3631_/Y vssd1 vssd1 vccd1 vccd1 _3657_/B sky130_fd_sc_hd__a21oi_2
X_6351_ _6401_/CLK _6351_/D vssd1 vssd1 vccd1 vccd1 _6351_/Q sky130_fd_sc_hd__dfxtp_1
X_3563_ _3563_/A _3563_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3564_/B sky130_fd_sc_hd__and3_1
X_5302_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5302_/X sky130_fd_sc_hd__or2_1
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3494_ _3525_/A _3494_/B _3685_/B vssd1 vssd1 vccd1 vccd1 _3494_/X sky130_fd_sc_hd__and3_1
XFILLER_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6282_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5233_ _5233_/A _5283_/A vssd1 vssd1 vccd1 vccd1 _5244_/B sky130_fd_sc_hd__and2_1
X_5164_ _5118_/A _5128_/B _5199_/B _5160_/Y vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__a31o_1
X_4115_ _4096_/B _4114_/X _5246_/A _3969_/X vssd1 vssd1 vccd1 vccd1 _4118_/C sky130_fd_sc_hd__o211ai_4
XFILLER_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5095_ _5095_/A _5168_/B vssd1 vssd1 vccd1 vccd1 _5137_/A sky130_fd_sc_hd__nand2_2
X_4046_ _4027_/X _4044_/X _3996_/X _4045_/Y vssd1 vssd1 vccd1 vccd1 _4050_/A sky130_fd_sc_hd__o211ai_2
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _5997_/A _5997_/B vssd1 vssd1 vccd1 vccd1 _6004_/B sky130_fd_sc_hd__xnor2_1
X_4948_ _4948_/A _4967_/B _4948_/C vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__and3_1
X_4879_ _4879_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _4879_/Y sky130_fd_sc_hd__nor2_1
X_6618_ _6618_/A _3313_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_6549_ _6549_/A _3233_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5920_ _6100_/A vssd1 vssd1 vccd1 vccd1 _6115_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ _5851_/A vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__buf_2
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4802_ _4802_/A _4802_/B _4813_/A _4802_/D vssd1 vssd1 vccd1 vccd1 _4813_/B sky130_fd_sc_hd__nand4_1
X_5782_ _6402_/Q _5782_/B vssd1 vssd1 vccd1 vccd1 _5784_/C sky130_fd_sc_hd__or2_1
X_4733_ _4733_/A vssd1 vssd1 vccd1 vccd1 _4734_/C sky130_fd_sc_hd__inv_2
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6403_ _6425_/CLK _6403_/D vssd1 vssd1 vccd1 vccd1 _6403_/Q sky130_fd_sc_hd__dfxtp_1
X_4664_ _4745_/A _4828_/A _4855_/B _4855_/C vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__nand4_2
X_4595_ _4594_/A _4594_/B _4594_/C vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__a21oi_1
X_3615_ _4677_/A _3716_/D _3650_/B vssd1 vssd1 vccd1 vccd1 _3615_/X sky130_fd_sc_hd__and3_1
X_3546_ _3546_/A _3546_/B vssd1 vssd1 vccd1 vccd1 _3588_/A sky130_fd_sc_hd__xor2_1
X_6334_ _6396_/CLK _6334_/D vssd1 vssd1 vccd1 vccd1 _6334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6265_ _6407_/Q _6268_/C vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__and2_1
X_3477_ _3477_/A _3477_/B vssd1 vssd1 vccd1 vccd1 _3479_/B sky130_fd_sc_hd__nor2_1
X_5216_ _5222_/A _5216_/B vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__xnor2_1
X_6196_ _6234_/A vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5147_ _5147_/A _5147_/B vssd1 vssd1 vccd1 vccd1 _5148_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _5079_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__or2_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4029_ _5492_/A vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ _4380_/A _4380_/B vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__xnor2_4
X_3400_ _4728_/A vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__buf_2
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3331_ _3333_/A vssd1 vssd1 vccd1 vccd1 _3331_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3266_/A vssd1 vssd1 vccd1 vccd1 _3262_/Y sky130_fd_sc_hd__inv_2
X_6050_ _6099_/A _6050_/B vssd1 vssd1 vccd1 vccd1 _6050_/Y sky130_fd_sc_hd__nand2_1
X_5001_ _5001_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5065_/B sky130_fd_sc_hd__xor2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5903_ _6426_/Q _6325_/Q vssd1 vssd1 vccd1 vccd1 _5903_/Y sky130_fd_sc_hd__nor2_1
X_5834_ _5828_/X _6410_/Q _5831_/X _5833_/Y vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__o31a_1
XFILLER_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5765_ _5916_/A vssd1 vssd1 vccd1 vccd1 _5765_/X sky130_fd_sc_hd__buf_2
X_4716_ _4769_/B vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__buf_2
X_5696_ _5785_/A _5717_/B _5695_/X vssd1 vssd1 vccd1 vccd1 _5696_/X sky130_fd_sc_hd__a21o_1
X_4647_ _4711_/D vssd1 vssd1 vccd1 vccd1 _4812_/B sky130_fd_sc_hd__clkbuf_2
X_4578_ _4578_/A _4379_/X vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__or2b_2
X_6317_ _6361_/CLK _6317_/D vssd1 vssd1 vccd1 vccd1 _6317_/Q sky130_fd_sc_hd__dfxtp_1
X_3529_ _3529_/A _3529_/B vssd1 vssd1 vccd1 vccd1 _3535_/A sky130_fd_sc_hd__or2_1
XFILLER_39_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6248_ _6398_/Q _6397_/Q _6400_/Q _6399_/Q vssd1 vssd1 vccd1 vccd1 _6248_/X sky130_fd_sc_hd__or4_1
X_6179_ _6367_/Q _6366_/Q _6178_/X _6324_/D vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__o31a_1
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3880_ _3891_/A _3891_/B _3879_/X vssd1 vssd1 vccd1 vccd1 _3882_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _5553_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _5550_/X sky130_fd_sc_hd__and2b_1
X_4501_ _4498_/Y _4484_/B _4500_/X vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__o21a_1
X_5481_ _5482_/B _5481_/B vssd1 vssd1 vccd1 vccd1 _5485_/B sky130_fd_sc_hd__xnor2_1
X_4432_ _4448_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4544_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4363_ _4363_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4374_/B sky130_fd_sc_hd__xnor2_2
X_3314_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3314_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4294_ _4294_/A _4294_/B vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6294_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3245_ _3247_/A vssd1 vssd1 vccd1 vccd1 _3245_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6041_/A vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ _5817_/A vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__clkbuf_1
X_5748_ _5748_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__xor2_2
XFILLER_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5679_ _5565_/X _5679_/B _5686_/A vssd1 vssd1 vccd1 vccd1 _5680_/B sky130_fd_sc_hd__and3b_1
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4981_ _4945_/B _4943_/X _4981_/S vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _5122_/A _4118_/B _3930_/C vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3863_ _4095_/A vssd1 vssd1 vccd1 vccd1 _5288_/A sky130_fd_sc_hd__clkbuf_2
X_6582_ _6582_/A _3272_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_5602_ _5602_/A _5602_/B vssd1 vssd1 vccd1 vccd1 _5605_/A sky130_fd_sc_hd__nand2_1
X_3794_ _3808_/B _3841_/A vssd1 vssd1 vccd1 vccd1 _3843_/A sky130_fd_sc_hd__nor2_1
X_5533_ _6317_/Q _5533_/B _5533_/C vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__and3_1
X_5464_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5465_/B sky130_fd_sc_hd__xnor2_1
X_4415_ _4415_/A _4415_/B vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__nor2_1
X_5395_ _5533_/B vssd1 vssd1 vccd1 vccd1 _5555_/D sky130_fd_sc_hd__buf_2
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4346_ _4345_/A _4368_/A _4368_/B _4366_/A _4366_/B vssd1 vssd1 vccd1 vccd1 _4350_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4277_ _5367_/A _4424_/B _4308_/B _4276_/A vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__a31o_1
X_3228_ _3229_/A vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6016_ _5756_/A _5982_/A _6014_/Y _6015_/X vssd1 vssd1 vccd1 vccd1 _6332_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4200_ _4200_/A _4200_/B _4246_/B vssd1 vssd1 vccd1 vccd1 _4201_/B sky130_fd_sc_hd__or3_1
X_5180_ _5257_/A _5180_/B vssd1 vssd1 vccd1 vccd1 _5182_/C sky130_fd_sc_hd__and2_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4131_ _4131_/A _4185_/A vssd1 vssd1 vccd1 vccd1 _4231_/A sky130_fd_sc_hd__xor2_1
X_4062_ _4104_/A _5237_/A _4373_/B _4212_/B vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__and4_1
XFILLER_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4964_ _5234_/A _5157_/B vssd1 vssd1 vccd1 vccd1 _5106_/B sky130_fd_sc_hd__or2b_2
X_3915_ _3915_/A _3915_/B _3992_/B _5697_/A vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__or4bb_1
X_4895_ _4895_/A _4895_/B _4895_/C _4895_/D vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__and4_1
X_6634_ _6634_/A _3338_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_3846_ _3812_/A _3846_/B vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__and2b_1
X_6565_ _6565_/A _3251_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
X_3777_ _3992_/B vssd1 vssd1 vccd1 vccd1 _4041_/B sky130_fd_sc_hd__buf_2
X_5516_ _5516_/A _5516_/B vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__xnor2_2
X_5447_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5447_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5378_ _5379_/B _5378_/B vssd1 vssd1 vccd1 vccd1 _5398_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4329_ _4329_/A _4329_/B vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3708_/A _3726_/A vssd1 vssd1 vccd1 vccd1 _3704_/A sky130_fd_sc_hd__xnor2_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4680_ _4684_/B _4680_/B vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__xnor2_1
X_3631_ _3593_/B _3630_/X _3660_/A vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__a21oi_1
X_3562_ _3563_/B _3563_/C _3563_/A vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__a21oi_1
X_6350_ _6401_/CLK _6350_/D vssd1 vssd1 vccd1 vccd1 _6350_/Q sky130_fd_sc_hd__dfxtp_1
X_5301_ _5301_/A _5301_/B vssd1 vssd1 vccd1 vccd1 _5341_/B sky130_fd_sc_hd__xor2_2
X_3493_ _3592_/C vssd1 vssd1 vccd1 vccd1 _3685_/B sky130_fd_sc_hd__clkbuf_2
X_6281_ _6413_/Q _6283_/C _6280_/Y vssd1 vssd1 vccd1 vccd1 _6413_/D sky130_fd_sc_hd__o21a_1
X_5232_ _5406_/A _5455_/B _5455_/C vssd1 vssd1 vccd1 vccd1 _5283_/A sky130_fd_sc_hd__and3_1
X_5163_ _5160_/Y _5163_/B vssd1 vssd1 vccd1 vccd1 _5199_/B sky130_fd_sc_hd__and2b_1
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4114_ _5248_/B _4221_/B _4114_/C vssd1 vssd1 vccd1 vccd1 _4114_/X sky130_fd_sc_hd__and3_1
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5094_ _5248_/D vssd1 vssd1 vccd1 vccd1 _5128_/B sky130_fd_sc_hd__buf_2
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4045_ _3996_/A _3996_/C _3996_/B vssd1 vssd1 vccd1 vccd1 _4045_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5996_ _4627_/A _5994_/X _5995_/Y vssd1 vssd1 vccd1 vccd1 _6329_/D sky130_fd_sc_hd__o21a_1
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4947_ _4978_/A _4978_/B _4978_/C vssd1 vssd1 vccd1 vccd1 _4979_/C sky130_fd_sc_hd__a21oi_2
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4878_ _4878_/A _4878_/B _4878_/C vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__nand3_2
X_6617_ _6617_/A _3311_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
X_3829_ _5281_/A vssd1 vssd1 vccd1 vccd1 _5198_/A sky130_fd_sc_hd__clkbuf_2
X_6548_ _6548_/A _3232_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6505__87 vssd1 vssd1 vccd1 vccd1 _6505__87/HI _6613_/A sky130_fd_sc_hd__conb_1
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _3364_/A _5750_/X _5849_/X _5748_/X vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5781_ _5829_/A _5746_/A _5780_/X _5868_/A vssd1 vssd1 vccd1 vccd1 _5782_/B sky130_fd_sc_hd__o2bb2a_1
X_4801_ _4830_/A _4830_/C _4800_/C vssd1 vssd1 vccd1 vccd1 _4802_/D sky130_fd_sc_hd__a21o_1
X_4732_ _4732_/A _4923_/B vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__xor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _4855_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3614_ _4855_/A vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__buf_2
X_6402_ _6425_/CLK _6402_/D vssd1 vssd1 vccd1 vccd1 _6402_/Q sky130_fd_sc_hd__dfxtp_1
X_4594_ _4594_/A _4594_/B _4594_/C vssd1 vssd1 vccd1 vccd1 _4614_/A sky130_fd_sc_hd__and3_1
X_3545_ _3547_/A _3547_/B _3548_/B vssd1 vssd1 vccd1 vccd1 _3553_/B sky130_fd_sc_hd__a21o_1
X_6333_ _6345_/CLK _6333_/D vssd1 vssd1 vccd1 vccd1 _6333_/Q sky130_fd_sc_hd__dfxtp_1
X_3476_ _3484_/B _3484_/A vssd1 vssd1 vccd1 vccd1 _3477_/B sky130_fd_sc_hd__and2b_1
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6264_ _6406_/Q _6260_/B _6263_/Y vssd1 vssd1 vccd1 vccd1 _6406_/D sky130_fd_sc_hd__o21a_1
XFILLER_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5215_ _5215_/A _5221_/A vssd1 vssd1 vccd1 vccd1 _5216_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6195_ _6195_/A vssd1 vssd1 vccd1 vccd1 _6381_/D sky130_fd_sc_hd__clkbuf_1
X_5146_ _5140_/A _5140_/B _5145_/X vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__a21bo_2
XFILLER_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5077_ _5136_/A _5101_/B vssd1 vssd1 vccd1 vccd1 _5079_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ _6316_/Q vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5979_ _5979_/A _5984_/A vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__or2_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3330_ _3333_/A vssd1 vssd1 vccd1 vccd1 _3330_/Y sky130_fd_sc_hd__inv_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A _5096_/B vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__and2_1
X_3261_ _3279_/A vssd1 vssd1 vccd1 vccd1 _3266_/A sky130_fd_sc_hd__buf_8
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5902_ _6426_/Q _6325_/Q vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__and2_1
X_5833_ _5765_/X _5825_/A _5832_/X _5807_/A vssd1 vssd1 vccd1 vccd1 _5833_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5764_ _6403_/Q vssd1 vssd1 vccd1 vccd1 _5783_/A sky130_fd_sc_hd__inv_2
X_4715_ _4715_/A _4715_/B vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__xnor2_1
X_5695_ _5695_/A _5695_/B vssd1 vssd1 vccd1 vccd1 _5695_/X sky130_fd_sc_hd__and2_1
X_4646_ _4769_/B _4646_/B vssd1 vssd1 vccd1 vccd1 _4711_/D sky130_fd_sc_hd__nor2_1
X_4577_ _4872_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _4905_/C sky130_fd_sc_hd__and2_2
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _6426_/CLK _6316_/D vssd1 vssd1 vccd1 vccd1 _6316_/Q sky130_fd_sc_hd__dfxtp_1
X_3528_ _4688_/B _3534_/D _3528_/C vssd1 vssd1 vccd1 vccd1 _3529_/B sky130_fd_sc_hd__and3_1
X_6496__78 vssd1 vssd1 vccd1 vccd1 _6496__78/HI _6604_/A sky130_fd_sc_hd__conb_1
X_3459_ _4677_/A vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6247_ _6394_/Q _6393_/Q _6396_/Q _6395_/Q vssd1 vssd1 vccd1 vccd1 _6247_/X sky130_fd_sc_hd__or4_1
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6178_ _6369_/Q _6368_/Q _6178_/C vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__or3_1
X_5129_ _5129_/A _5129_/B vssd1 vssd1 vccd1 vccd1 _5152_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5480_ _5494_/A _5494_/B _5479_/X vssd1 vssd1 vccd1 vccd1 _5481_/B sky130_fd_sc_hd__o21ba_1
X_4500_ _3887_/B _3849_/Y _3853_/B _3887_/A _4499_/Y vssd1 vssd1 vccd1 vccd1 _4500_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4431_ _4431_/A _4445_/A vssd1 vssd1 vccd1 vccd1 _4448_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4362_ _5545_/A _4391_/B _4391_/C vssd1 vssd1 vccd1 vccd1 _4364_/B sky130_fd_sc_hd__and3_1
X_4293_ _4463_/B _4293_/B vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__xnor2_4
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3313_/Y sky130_fd_sc_hd__inv_2
X_6101_ _6104_/A _6032_/X _6097_/X _6099_/Y _6100_/X vssd1 vssd1 vccd1 vccd1 _6345_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3244_ _3247_/A vssd1 vssd1 vccd1 vccd1 _3244_/Y sky130_fd_sc_hd__inv_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6041_/A vssd1 vssd1 vccd1 vccd1 _6032_/X sky130_fd_sc_hd__clkbuf_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5816_ _5871_/B vssd1 vssd1 vccd1 vccd1 _6104_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5747_ _5803_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _5684_/A vssd1 vssd1 vccd1 vccd1 _5842_/A sky130_fd_sc_hd__buf_2
X_4629_ _4629_/A _4629_/B vssd1 vssd1 vccd1 vccd1 _4630_/C sky130_fd_sc_hd__or2_1
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _4980_/A _4946_/B vssd1 vssd1 vccd1 vccd1 _4983_/C sky130_fd_sc_hd__or2b_1
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _3931_/A vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3862_ _5322_/A vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6581_ _6581_/A _3271_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_32_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5601_ _5601_/A _5050_/B vssd1 vssd1 vccd1 vccd1 _5602_/B sky130_fd_sc_hd__or2b_1
X_3793_ _5211_/A _3858_/B vssd1 vssd1 vccd1 vccd1 _3841_/A sky130_fd_sc_hd__nand2_1
X_5532_ _5532_/A _5532_/B vssd1 vssd1 vccd1 vccd1 _5533_/C sky130_fd_sc_hd__xnor2_1
X_5463_ _5466_/A _5466_/B _5462_/A vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__a21o_1
X_5394_ _5394_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__nand2_1
X_4414_ _5458_/A _4188_/X _4387_/C vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__a21oi_1
X_4345_ _4345_/A _4345_/B vssd1 vssd1 vccd1 vccd1 _4366_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _4276_/A _4276_/B vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__nor2_1
X_6466__48 vssd1 vssd1 vccd1 vccd1 _6466__48/HI _6571_/A sky130_fd_sc_hd__conb_1
X_3227_ _3229_/A vssd1 vssd1 vccd1 vccd1 _3227_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6015_ _6115_/B vssd1 vssd1 vccd1 vccd1 _6015_/X sky130_fd_sc_hd__buf_2
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6480__62 vssd1 vssd1 vccd1 vccd1 _6480__62/HI _6588_/A sky130_fd_sc_hd__conb_1
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4130_ _5159_/A _4109_/B _4109_/C vssd1 vssd1 vccd1 vccd1 _4144_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4061_ _4104_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _4963_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _5157_/B sky130_fd_sc_hd__xnor2_4
X_3914_ _5068_/A vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__buf_2
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6633_ _6633_/A _3340_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4894_ _4909_/A _4909_/B _4909_/C vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3845_ _3855_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3887_/A sky130_fd_sc_hd__or2_2
X_6564_ _6564_/A _3342_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
X_3776_ _3385_/Y _3442_/A _3445_/A _3775_/X vssd1 vssd1 vccd1 vccd1 _3992_/B sky130_fd_sc_hd__o22a_4
X_5515_ _5511_/Y _5514_/X _4373_/A _5317_/B vssd1 vssd1 vccd1 vccd1 _5530_/A sky130_fd_sc_hd__o211ai_4
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5446_ _5438_/X _5439_/Y _5468_/B _5445_/B _5445_/A vssd1 vssd1 vccd1 vccd1 _5464_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5377_ _5400_/A _5400_/B _5376_/X vssd1 vssd1 vccd1 vccd1 _5378_/B sky130_fd_sc_hd__o21ba_1
XFILLER_101_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4328_ _4321_/A _4327_/X _4349_/A vssd1 vssd1 vccd1 vccd1 _4328_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4259_ _5386_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4266_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3630_ _3672_/A _3592_/C _4694_/B _3699_/A vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__a22o_1
X_3561_ _3561_/A _3561_/B vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__nand2_1
X_5300_ _5300_/A _5305_/B vssd1 vssd1 vccd1 vccd1 _5301_/B sky130_fd_sc_hd__xnor2_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3492_ _3502_/B vssd1 vssd1 vccd1 vccd1 _3544_/A sky130_fd_sc_hd__inv_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6280_ _6280_/A _6280_/B vssd1 vssd1 vccd1 vccd1 _6280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5231_ _5231_/A _5231_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5455_/C sky130_fd_sc_hd__or3_2
XFILLER_96_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5162_ _5102_/A _5288_/B _5240_/B _5282_/A vssd1 vssd1 vccd1 vccd1 _5163_/B sky130_fd_sc_hd__a22o_1
X_6436__18 vssd1 vssd1 vccd1 vccd1 _6436__18/HI _6541_/A sky130_fd_sc_hd__conb_1
X_4113_ _4113_/A _4113_/B _4113_/C vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__or3_4
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5093_ _5392_/B vssd1 vssd1 vccd1 vccd1 _5248_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4044_ _4027_/X _4047_/B _4044_/C _4044_/D vssd1 vssd1 vccd1 vccd1 _4044_/X sky130_fd_sc_hd__and4b_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5995_ _4627_/A _5994_/X _6299_/A vssd1 vssd1 vccd1 vccd1 _5995_/Y sky130_fd_sc_hd__a21oi_1
X_4946_ _4946_/A _4946_/B vssd1 vssd1 vccd1 vccd1 _4978_/C sky130_fd_sc_hd__xnor2_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4877_ _4885_/A _4885_/B vssd1 vssd1 vccd1 vccd1 _4878_/C sky130_fd_sc_hd__nor2_1
X_3828_ _4212_/A vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__clkbuf_2
X_6616_ _6616_/A _3308_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_6547_ _6547_/A _3231_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3759_ _3759_/A _3759_/B _3759_/C vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__and3_1
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5429_ _5560_/A _5288_/B _5428_/C vssd1 vssd1 vccd1 vccd1 _5430_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6450__32 vssd1 vssd1 vccd1 vccd1 _6450__32/HI _6555_/A sky130_fd_sc_hd__conb_1
XFILLER_70_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4800_ _4800_/A _4830_/C _4800_/C vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__nand3_1
XFILLER_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5780_ _5823_/B _5775_/Y _5779_/Y _5751_/Y vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4728_/A _4834_/B _4712_/X _4713_/A vssd1 vssd1 vccd1 vccd1 _4923_/B sky130_fd_sc_hd__a31o_1
X_4662_ _4660_/B _4648_/B _3628_/C vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__o21ai_1
X_6401_ _6401_/CLK _6401_/D vssd1 vssd1 vccd1 vccd1 _6401_/Q sky130_fd_sc_hd__dfxtp_1
X_3613_ _3627_/A _3627_/B _3610_/X vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__a21bo_1
X_4593_ _4542_/X _4549_/X _4591_/X _4592_/X vssd1 vssd1 vccd1 vccd1 _4593_/X sky130_fd_sc_hd__a31o_1
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3544_ _3544_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3548_/B sky130_fd_sc_hd__and2_1
X_6332_ _6361_/CLK _6332_/D vssd1 vssd1 vccd1 vccd1 _6332_/Q sky130_fd_sc_hd__dfxtp_1
X_3475_ _3480_/A _3475_/B vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__nand2_1
X_6263_ _6280_/A _6268_/C vssd1 vssd1 vccd1 vccd1 _6263_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5214_ _5214_/A _5214_/B vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6194_ _6380_/Q _6194_/B vssd1 vssd1 vccd1 vccd1 _6195_/A sky130_fd_sc_hd__and2_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5145_ _5145_/A _5135_/B vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__or2b_1
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5076_ _5081_/B _5076_/B vssd1 vssd1 vccd1 vccd1 _5147_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4027_ _4027_/A _4027_/B _4027_/C vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__and3_1
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5978_ _5978_/A _5984_/A vssd1 vssd1 vccd1 vccd1 _5978_/X sky130_fd_sc_hd__and2_1
XFILLER_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4929_/A _4929_/B vssd1 vssd1 vccd1 vccd1 _4931_/C sky130_fd_sc_hd__xnor2_1
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3260_/A vssd1 vssd1 vccd1 vccd1 _3260_/Y sky130_fd_sc_hd__inv_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5890_/X _5898_/X _5900_/Y vssd1 vssd1 vccd1 vccd1 _6578_/A sky130_fd_sc_hd__a21oi_2
XFILLER_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5832_ _5818_/X _5769_/Y _5820_/X _5767_/X vssd1 vssd1 vccd1 vccd1 _5832_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5763_ _6404_/Q _5793_/B vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__and2_1
X_4714_ _4714_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4715_/B sky130_fd_sc_hd__xnor2_1
X_5694_ _5695_/A _5695_/B vssd1 vssd1 vccd1 vccd1 _5717_/B sky130_fd_sc_hd__xor2_1
X_4645_ _6074_/A _4751_/C _4643_/C vssd1 vssd1 vccd1 vccd1 _4646_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4576_ _4596_/C _4580_/B vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3527_ _4688_/B _3534_/D _3528_/C vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__a21oi_1
X_6315_ _6315_/A vssd1 vssd1 vccd1 vccd1 _6426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3458_ _3395_/A _3494_/B _3466_/B _4651_/A vssd1 vssd1 vccd1 vccd1 _3462_/A sky130_fd_sc_hd__a22o_1
X_6246_ _6393_/Q _6396_/Q _6246_/C vssd1 vssd1 vccd1 vccd1 _6246_/X sky130_fd_sc_hd__and3_1
XFILLER_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3389_ _3525_/A vssd1 vssd1 vccd1 vccd1 _6010_/A sky130_fd_sc_hd__inv_2
X_6177_ _6371_/Q _6370_/Q _6373_/Q _6372_/Q vssd1 vssd1 vccd1 vccd1 _6178_/C sky130_fd_sc_hd__or4_1
X_5128_ _5136_/A _5128_/B vssd1 vssd1 vccd1 vccd1 _5129_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5290_/B vssd1 vssd1 vccd1 vccd1 _5353_/B sky130_fd_sc_hd__buf_2
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ _4433_/A _4433_/B vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4361_ _5518_/A vssd1 vssd1 vccd1 vccd1 _5545_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6100_ _6100_/A vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__clkbuf_4
X_4292_ _4292_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4293_/B sky130_fd_sc_hd__nor2_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3312_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3247_/A vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__inv_2
X_6031_ _6027_/X _6028_/Y _6029_/X _6030_/X vssd1 vssd1 vccd1 vccd1 _6041_/A sky130_fd_sc_hd__o22a_2
XFILLER_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5815_ _5815_/A vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5746_ _5746_/A vssd1 vssd1 vccd1 vccd1 _5746_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5677_ _5950_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _5677_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4628_ _4710_/A vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4559_ _4567_/A _4559_/B vssd1 vssd1 vccd1 vccd1 _4560_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6229_ _6229_/A vssd1 vssd1 vccd1 vccd1 _6393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _5096_/A _3931_/A _3930_/C vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__and3_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3861_ _5456_/A vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__clkbuf_2
X_3792_ _3903_/B vssd1 vssd1 vccd1 vccd1 _3858_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6580_ _6580_/A _3270_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
X_5600_ _5600_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5803_/A sky130_fd_sc_hd__xnor2_4
XFILLER_31_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5531_ _5531_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__xnor2_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5462_ _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _5466_/B sky130_fd_sc_hd__nor2_1
X_5393_ _5392_/A _5392_/B _5392_/C vssd1 vssd1 vccd1 vccd1 _5394_/B sky130_fd_sc_hd__a21o_1
X_4413_ _4413_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4344_ _4368_/A _4368_/B vssd1 vssd1 vccd1 vccd1 _4345_/B sky130_fd_sc_hd__or2_1
XFILLER_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4275_ _5441_/A _4336_/A _5466_/A vssd1 vssd1 vccd1 vccd1 _4276_/B sky130_fd_sc_hd__a21oi_1
X_6014_ _6014_/A _6014_/B vssd1 vssd1 vccd1 vccd1 _6014_/Y sky130_fd_sc_hd__nand2_1
X_3226_ _3229_/A vssd1 vssd1 vccd1 vccd1 _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5729_ _5729_/A _5729_/B _5728_/X vssd1 vssd1 vccd1 vccd1 _5729_/X sky130_fd_sc_hd__or3b_1
XFILLER_117_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4060_ _4213_/D vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _5193_/A _5193_/B _5230_/A vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__o21bai_4
X_3913_ _3974_/A vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__clkbuf_2
X_4893_ _4907_/A _4907_/B vssd1 vssd1 vccd1 vccd1 _4909_/C sky130_fd_sc_hd__and2b_1
X_6632_ _6632_/A _3331_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_3844_ _3844_/A _3844_/B vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6563_ _6563_/A _3250_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
X_3775_ _3791_/A _3791_/B vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5514_ _5514_/A _5514_/B _5519_/A vssd1 vssd1 vccd1 vccd1 _5514_/X sky130_fd_sc_hd__and3_1
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5445_ _5445_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5468_/B sky130_fd_sc_hd__xnor2_2
XFILLER_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5376_ _5375_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__and2b_1
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4327_ _4327_/A _4327_/B vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__and2_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4258_ _5691_/A _4256_/Y _4297_/A _4257_/X vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__o31ai_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ input1/X vssd1 vssd1 vccd1 vccd1 _3334_/A sky130_fd_sc_hd__clkbuf_4
X_4189_ _4272_/A _4424_/B _4183_/X vssd1 vssd1 vccd1 vccd1 _4189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3560_ _3560_/A _3560_/B vssd1 vssd1 vccd1 vccd1 _3561_/B sky130_fd_sc_hd__nand2_1
X_3491_ _3646_/A _3699_/A _3592_/D _4643_/C vssd1 vssd1 vccd1 vccd1 _3502_/B sky130_fd_sc_hd__and4_2
X_5230_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5455_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5161_ _5460_/B vssd1 vssd1 vccd1 vccd1 _5240_/B sky130_fd_sc_hd__buf_2
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4112_ _4149_/A _4148_/B _4111_/X vssd1 vssd1 vccd1 vccd1 _4113_/C sky130_fd_sc_hd__a21oi_1
X_5092_ _5092_/A _5092_/B vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4043_ _4027_/A _4027_/B _4027_/C vssd1 vssd1 vccd1 vccd1 _4044_/D sky130_fd_sc_hd__a21o_1
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _6001_/S _5994_/B _5994_/C vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__and3_1
X_4945_ _4943_/X _4945_/B vssd1 vssd1 vccd1 vccd1 _4946_/B sky130_fd_sc_hd__and2b_1
XFILLER_33_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4876_ _4879_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__xnor2_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3827_ _5407_/A vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6615_ _6615_/A _3306_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_6546_ _6546_/A _3229_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_3758_ _4101_/B _4101_/C _4101_/A vssd1 vssd1 vccd1 vccd1 _3758_/X sky130_fd_sc_hd__a21bo_1
X_3689_ _3708_/A _3689_/B vssd1 vssd1 vccd1 vccd1 _3691_/B sky130_fd_sc_hd__xnor2_1
X_5428_ _5428_/A _5428_/B _5428_/C vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__and3_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5359_ _5359_/A _5359_/B vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__xor2_2
XFILLER_114_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4927_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__or2_1
X_4661_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3612_ _3612_/A _3716_/C vssd1 vssd1 vccd1 vccd1 _3627_/B sky130_fd_sc_hd__nand2_2
X_6400_ _6401_/CLK _6400_/D vssd1 vssd1 vccd1 vccd1 _6400_/Q sky130_fd_sc_hd__dfxtp_1
X_4592_ _4601_/B _4592_/B _4592_/C vssd1 vssd1 vccd1 vccd1 _4592_/X sky130_fd_sc_hd__and3_1
X_6331_ _6345_/CLK _6331_/D vssd1 vssd1 vccd1 vccd1 _6331_/Q sky130_fd_sc_hd__dfxtp_1
X_3543_ _4800_/A _3406_/B _3430_/B _4895_/A vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__a22o_1
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3474_ _4710_/A _3509_/B _3461_/A vssd1 vssd1 vccd1 vccd1 _3475_/B sky130_fd_sc_hd__a21o_1
X_6262_ _6406_/Q _6405_/Q _6262_/C vssd1 vssd1 vccd1 vccd1 _6268_/C sky130_fd_sc_hd__and3_1
X_5213_ _4581_/A _5299_/B _5205_/B _5212_/Y vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__a31o_1
X_6193_ _6193_/A vssd1 vssd1 vccd1 vccd1 _6380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5144_ _5144_/A _5144_/B vssd1 vssd1 vccd1 vccd1 _5591_/A sky130_fd_sc_hd__or2_2
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5075_ _5075_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _5076_/B sky130_fd_sc_hd__xor2_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4026_ _4024_/A _4024_/B _4075_/A vssd1 vssd1 vccd1 vccd1 _4027_/C sky130_fd_sc_hd__a21bo_1
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5977_ _5968_/X _5970_/X _5971_/X _5969_/Y vssd1 vssd1 vccd1 vccd1 _5984_/A sky130_fd_sc_hd__o22a_1
X_4928_ _4928_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4929_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4859_/A _4878_/A vssd1 vssd1 vccd1 vccd1 _4861_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6510__92 vssd1 vssd1 vccd1 vccd1 _6510__92/HI _6618_/A sky130_fd_sc_hd__conb_1
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5900_ _5893_/Y _5892_/X _5896_/Y _5899_/Y vssd1 vssd1 vccd1 vccd1 _5900_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5831_ _5918_/A _5825_/A _5830_/X _5743_/A vssd1 vssd1 vccd1 vccd1 _5831_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5762_ _5771_/A _5760_/X _5746_/A _5926_/A vssd1 vssd1 vccd1 vccd1 _5793_/B sky130_fd_sc_hd__a22oi_2
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4713_ _4713_/A _4712_/X vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__or2b_1
X_5693_ _5693_/A _5693_/B vssd1 vssd1 vccd1 vccd1 _5695_/B sky130_fd_sc_hd__xnor2_1
X_4644_ _6342_/Q vssd1 vssd1 vccd1 vccd1 _6074_/A sky130_fd_sc_hd__buf_2
XFILLER_116_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4575_ _4575_/A _4575_/B vssd1 vssd1 vccd1 vccd1 _4580_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3526_ _3546_/A _3546_/B _3523_/X vssd1 vssd1 vccd1 vccd1 _3528_/C sky130_fd_sc_hd__o21a_1
X_6314_ _6356_/Q _6314_/B vssd1 vssd1 vccd1 vccd1 _6315_/A sky130_fd_sc_hd__and2_1
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6245_ _6398_/Q _6397_/Q _6400_/Q _6399_/Q vssd1 vssd1 vccd1 vccd1 _6246_/C sky130_fd_sc_hd__and4_1
XFILLER_103_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3457_ _3699_/C vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__clkbuf_2
X_3388_ _3525_/A _3430_/B vssd1 vssd1 vccd1 vccd1 _3406_/C sky130_fd_sc_hd__and2_1
X_6176_ _6367_/Q _6366_/Q _6369_/Q _6368_/Q vssd1 vssd1 vccd1 vccd1 _6176_/X sky130_fd_sc_hd__and4_1
X_5127_ _5127_/A _5127_/B vssd1 vssd1 vccd1 vccd1 _5152_/A sky130_fd_sc_hd__xor2_1
X_5058_ _5290_/B vssd1 vssd1 vccd1 vccd1 _5297_/B sky130_fd_sc_hd__clkbuf_4
X_4009_ _4009_/A _4009_/B vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6487__69 vssd1 vssd1 vccd1 vccd1 _6487__69/HI _6595_/A sky130_fd_sc_hd__conb_1
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4360_ _4369_/A _4370_/B _4369_/B vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__o21ba_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3311_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4291_ _4294_/A _4294_/B vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__and2b_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3248_/A vssd1 vssd1 vccd1 vccd1 _3247_/A sky130_fd_sc_hd__buf_12
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6030_ _6392_/Q _6401_/Q vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__and2b_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5814_ _6409_/Q _5744_/X _5754_/X _5811_/X _6299_/A vssd1 vssd1 vccd1 vccd1 _6580_/A
+ sky130_fd_sc_hd__a221oi_4
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5745_ _5745_/A _5745_/B vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__or2_1
X_5676_ _5851_/A _5677_/B _5675_/X vssd1 vssd1 vccd1 vccd1 _5676_/X sky130_fd_sc_hd__a21o_1
X_4627_ _4627_/A _5985_/A vssd1 vssd1 vccd1 vccd1 _5756_/C sky130_fd_sc_hd__or2_1
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4558_ _5691_/A _4558_/B vssd1 vssd1 vccd1 vccd1 _4565_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3509_ _4629_/B _3509_/B vssd1 vssd1 vccd1 vccd1 _3515_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4489_ _4488_/B _4488_/C _4488_/A vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6228_ _6228_/A input6/X vssd1 vssd1 vccd1 vccd1 _6229_/A sky130_fd_sc_hd__and2_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6159_ _6159_/A vssd1 vssd1 vccd1 vccd1 _6366_/D sky130_fd_sc_hd__clkbuf_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3860_ _5487_/A vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__clkbuf_2
X_3791_ _3791_/A _3791_/B vssd1 vssd1 vccd1 vccd1 _3903_/B sky130_fd_sc_hd__xnor2_4
XFILLER_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5530_ _5530_/A _5530_/B vssd1 vssd1 vccd1 vccd1 _5568_/A sky130_fd_sc_hd__xnor2_2
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5461_ _5428_/A _5460_/B _5460_/C vssd1 vssd1 vccd1 vccd1 _5462_/B sky130_fd_sc_hd__a21oi_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4412_ _5492_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4413_/B sky130_fd_sc_hd__nand2_1
X_5392_ _5392_/A _5392_/B _5392_/C vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__nand3_1
X_4343_ _4347_/C _4343_/B vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__xor2_4
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4274_ _4274_/A _4573_/B vssd1 vssd1 vccd1 vccd1 _5466_/A sky130_fd_sc_hd__nor2_2
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3225_ _3229_/A vssd1 vssd1 vccd1 vccd1 _3225_/Y sky130_fd_sc_hd__inv_2
X_6013_ _6013_/A _6013_/B vssd1 vssd1 vccd1 vccd1 _6014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3989_ _5246_/A vssd1 vssd1 vccd1 vccd1 _5168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5728_ _5672_/Y _5676_/X _5727_/Y _5668_/X vssd1 vssd1 vccd1 vccd1 _5728_/X sky130_fd_sc_hd__o211a_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5659_ _5659_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5659_/X sky130_fd_sc_hd__or2_1
XFILLER_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6457__39 vssd1 vssd1 vccd1 vccd1 _6457__39/HI _6562_/A sky130_fd_sc_hd__conb_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6471__53 vssd1 vssd1 vccd1 vccd1 _6471__53/HI _6576_/A sky130_fd_sc_hd__conb_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _5231_/A _5231_/B _5231_/C vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__o21ai_1
X_3912_ _5248_/B vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4892_ _4900_/A _4899_/B _4899_/A vssd1 vssd1 vccd1 vccd1 _4907_/B sky130_fd_sc_hd__a21bo_1
X_6631_ _6631_/A _3330_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_3843_ _3843_/A _3843_/B _3843_/C vssd1 vssd1 vccd1 vccd1 _3844_/B sky130_fd_sc_hd__or3_1
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3774_ _3483_/X _3788_/B _3787_/A vssd1 vssd1 vccd1 vccd1 _3791_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6562_ _6562_/A _3249_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_5513_ _5511_/A _5532_/A _5512_/X vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__o21a_1
X_5444_ _5317_/A _5555_/D _5470_/B _5443_/A vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__a31oi_4
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5375_ _5375_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5400_/B sky130_fd_sc_hd__xor2_2
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4326_ _4326_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _4459_/B sky130_fd_sc_hd__xor2_4
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4257_ _5456_/A _4391_/B _4391_/C _4298_/B _5471_/A vssd1 vssd1 vccd1 vccd1 _4257_/X
+ sky130_fd_sc_hd__a32o_1
X_4188_ _4424_/B vssd1 vssd1 vccd1 vccd1 _4188_/X sky130_fd_sc_hd__buf_2
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3490_ _6327_/Q vssd1 vssd1 vccd1 vccd1 _3699_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ _5160_/A _5195_/A vssd1 vssd1 vccd1 vccd1 _5160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4111_ _4110_/B _4144_/A _4110_/A vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5091_ _5091_/A _5091_/B vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__nor2_2
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4042_ _5214_/A _4041_/B _4047_/A _4041_/D vssd1 vssd1 vccd1 vccd1 _4044_/C sky130_fd_sc_hd__a22o_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5993_ _5985_/A _5978_/A _5981_/A _5992_/X vssd1 vssd1 vccd1 vccd1 _5994_/C sky130_fd_sc_hd__o31ai_1
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ _4623_/A _4716_/X _4924_/B _3466_/A vssd1 vssd1 vccd1 vccd1 _4945_/B sky130_fd_sc_hd__a22o_1
X_4875_ _4875_/A _4875_/B vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__xor2_2
X_3826_ _5471_/A vssd1 vssd1 vccd1 vccd1 _5407_/A sky130_fd_sc_hd__buf_2
X_6614_ _6614_/A _3303_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_6545_ _6545_/A _3228_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_3757_ _3757_/A _3757_/B _3757_/C vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__nand3_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3688_ _4673_/B _3716_/D vssd1 vssd1 vccd1 vccd1 _3708_/A sky130_fd_sc_hd__nand2_1
X_5427_ _5390_/B _5475_/A _5467_/B _5426_/X vssd1 vssd1 vccd1 vccd1 _5428_/C sky130_fd_sc_hd__a22o_1
X_5358_ _5358_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _4404_/A _6321_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _5441_/C sky130_fd_sc_hd__and3_1
X_5289_ _5289_/A _5289_/B vssd1 vssd1 vccd1 vccd1 _5297_/C sky130_fd_sc_hd__xor2_2
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6441__23 vssd1 vssd1 vccd1 vccd1 _6441__23/HI _6546_/A sky130_fd_sc_hd__conb_1
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _6340_/Q _4660_/B _4660_/C vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__or3_2
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ _5997_/A _3608_/Y _3610_/X vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__o21a_1
X_4591_ _4549_/A _4549_/B _4557_/X _4590_/X vssd1 vssd1 vccd1 vccd1 _4591_/X sky130_fd_sc_hd__a22o_1
X_6330_ _6345_/CLK _6330_/D vssd1 vssd1 vccd1 vccd1 _6330_/Q sky130_fd_sc_hd__dfxtp_1
X_3542_ _3699_/A vssd1 vssd1 vccd1 vccd1 _4895_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3473_ _4805_/A _3473_/B _3473_/C vssd1 vssd1 vccd1 vccd1 _3480_/A sky130_fd_sc_hd__or3_2
X_6261_ _6405_/Q _6262_/C _6260_/Y vssd1 vssd1 vccd1 vccd1 _6405_/D sky130_fd_sc_hd__o21a_1
X_5212_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6192_ _6379_/Q _6194_/B vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__and2_1
X_5143_ _5151_/A _5151_/B _5142_/X vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__a21bo_2
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5074_ _5074_/A _5074_/B vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__nor2_1
X_4025_ _4037_/A _4025_/B _4025_/C vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__nand3_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5976_ _5981_/A _5982_/A _5975_/Y vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__a21oi_2
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4927_ _4927_/A _4927_/B vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _4859_/A _4858_/B _4858_/C vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__nand3_1
X_3809_ _5030_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _3810_/A sky130_fd_sc_hd__nand2_1
X_4789_ _4789_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5830_ _5775_/Y _5868_/C _5779_/Y _3364_/A vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5761_/A vssd1 vssd1 vccd1 vccd1 _5926_/A sky130_fd_sc_hd__buf_2
X_4712_ _4711_/A _4872_/B _4728_/B _4629_/B vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__a22o_1
X_5692_ _5692_/A _5699_/A vssd1 vssd1 vccd1 vccd1 _5693_/B sky130_fd_sc_hd__nor2_1
X_4643_ _6342_/Q _4751_/C _4643_/C vssd1 vssd1 vccd1 vccd1 _4769_/B sky130_fd_sc_hd__nor3_4
XFILLER_116_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4574_ _5712_/A _4436_/B _5560_/C vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3525_ _3525_/A _3718_/D vssd1 vssd1 vccd1 vccd1 _3546_/B sky130_fd_sc_hd__and2_1
X_6313_ _6425_/Q _6310_/B _6312_/Y vssd1 vssd1 vccd1 vccd1 _6425_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6400_/D sky130_fd_sc_hd__clkbuf_1
X_3456_ _3566_/A vssd1 vssd1 vccd1 vccd1 _3699_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3387_ _4756_/A vssd1 vssd1 vccd1 vccd1 _3525_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6175_ _6371_/Q _6370_/Q _6373_/Q _6372_/Q vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__and4_1
X_5126_ _5126_/A _5126_/B vssd1 vssd1 vccd1 vccd1 _5127_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5057_ _5057_/A _5057_/B vssd1 vssd1 vccd1 vccd1 _5290_/B sky130_fd_sc_hd__xnor2_4
X_4008_ _5102_/A _4008_/B vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5959_ _3354_/X _5933_/B _5956_/X _5957_/Y _6282_/A vssd1 vssd1 vccd1 vccd1 _5959_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3310_ _3310_/A vssd1 vssd1 vccd1 vccd1 _3315_/A sky130_fd_sc_hd__buf_12
X_4290_ _4290_/A _4290_/B vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__xnor2_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3241_/A vssd1 vssd1 vccd1 vccd1 _3241_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5813_ _6310_/A vssd1 vssd1 vccd1 vccd1 _6299_/A sky130_fd_sc_hd__buf_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5744_ _4635_/X _5742_/Y _5743_/X _4274_/A vssd1 vssd1 vccd1 vccd1 _5744_/X sky130_fd_sc_hd__a2bb2o_1
X_5675_ _5674_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__and2b_1
X_4626_ _4682_/A vssd1 vssd1 vccd1 vccd1 _5985_/A sky130_fd_sc_hd__clkbuf_2
X_4557_ _4557_/A _4557_/B vssd1 vssd1 vccd1 vccd1 _4557_/X sky130_fd_sc_hd__or2_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3508_ _4711_/B vssd1 vssd1 vccd1 vccd1 _4629_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4488_ _4488_/A _4488_/B _4488_/C vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__and3_1
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3439_ _4623_/A _3509_/B _3446_/C vssd1 vssd1 vccd1 vccd1 _3447_/A sky130_fd_sc_hd__a21oi_1
X_6227_ _6385_/Q _6386_/Q _6100_/X _6223_/X _6226_/X vssd1 vssd1 vccd1 vccd1 _6392_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6158_ _6228_/A input3/X vssd1 vssd1 vccd1 vccd1 _6159_/A sky130_fd_sc_hd__and2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5109_ _5110_/A _5160_/A vssd1 vssd1 vccd1 vccd1 _5155_/B sky130_fd_sc_hd__xor2_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6097_/A _6089_/B vssd1 vssd1 vccd1 vccd1 _6092_/A sky130_fd_sc_hd__and2_1
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3790_ _5030_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3808_/B sky130_fd_sc_hd__nand2_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5460_ _5555_/C _5460_/B _5460_/C vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__and3_1
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4411_ _4411_/A _4411_/B vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__xnor2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _5401_/A _5401_/B _5390_/Y vssd1 vssd1 vccd1 vccd1 _5392_/C sky130_fd_sc_hd__o21ai_1
X_4342_ _4373_/A _4342_/B vssd1 vssd1 vccd1 vccd1 _4343_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4273_ _6323_/Q vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__clkinv_4
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3224_ _3248_/A vssd1 vssd1 vccd1 vccd1 _3229_/A sky130_fd_sc_hd__buf_12
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6012_ _4629_/A _5992_/X _6011_/X vssd1 vssd1 vccd1 vccd1 _6013_/B sky130_fd_sc_hd__o21a_1
.ends

