* NGSPICE file created from wrapped_hsv_mixer.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt wrapped_hsv_mixer active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5469__C _5469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6286__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5766__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3988_ _3993_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _3994_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5485__B _5485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _5727_/A _5792_/A vssd1 vssd1 vccd1 vccd1 _5727_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3286__A _3288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5658_ _5659_/A _5659_/B _5657_/Y vssd1 vssd1 vccd1 vccd1 _5658_/Y sky130_fd_sc_hd__o21ai_1
X_4609_ _4613_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4609_/Y sky130_fd_sc_hd__nor2_1
X_5589_ _5589_/A _5589_/B vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__xnor2_2
XFILLER_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3196__A _3321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4960_/A _5000_/B vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3425__A2 _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3911_ _3911_/A _3923_/C vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__xor2_1
X_4891_ _4891_/A _4908_/A vssd1 vssd1 vccd1 vccd1 _4910_/C sky130_fd_sc_hd__nand2_1
X_3842_ _5037_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _3961_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6561_ _6561_/A _3275_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_3773_ _3773_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3774_/B sky130_fd_sc_hd__nor2_1
X_5512_ _5512_/A _5512_/B _5365_/X vssd1 vssd1 vccd1 vccd1 _5514_/B sky130_fd_sc_hd__or3b_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6492_ _6492_/A _3193_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_5443_ _5445_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5447_/A sky130_fd_sc_hd__or2b_1
X_5374_ _5380_/A _5380_/B _5373_/X vssd1 vssd1 vccd1 vccd1 _5376_/B sky130_fd_sc_hd__a21bo_1
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4325_ _4306_/A _4323_/Y _4324_/Y vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__o21ai_4
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4256_ _4257_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__xor2_4
XFILLER_101_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3207_ _3208_/A vssd1 vssd1 vccd1 vccd1 _3207_/Y sky130_fd_sc_hd__inv_2
X_4187_ _4187_/A _4187_/B vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__xor2_2
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4665__A _4769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_475 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6301__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_58 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5090_ _5231_/D vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__clkbuf_2
X_4110_ _3614_/Y _4110_/B vssd1 vssd1 vccd1 vccd1 _4110_/X sky130_fd_sc_hd__and2b_1
XFILLER_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4041_ _4042_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _4041_/X sky130_fd_sc_hd__and2_1
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ _5982_/X _5984_/X _5985_/X _5983_/Y vssd1 vssd1 vccd1 vccd1 _6000_/B sky130_fd_sc_hd__o22a_1
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4943_ _4923_/A _4923_/B _4705_/A vssd1 vssd1 vccd1 vccd1 _4944_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4874_ _4860_/B _4862_/X _4873_/A _4910_/A vssd1 vssd1 vccd1 vccd1 _5125_/B sky130_fd_sc_hd__o211ai_2
X_3825_ _3825_/A _3825_/B vssd1 vssd1 vccd1 vccd1 _3826_/B sky130_fd_sc_hd__xnor2_4
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3756_ _4929_/A _4168_/B _3754_/B _3755_/X vssd1 vssd1 vccd1 vccd1 _3793_/A sky130_fd_sc_hd__a31o_1
X_6544_ _6544_/A _3317_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3687_ _3687_/A _3693_/A vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__nand2_1
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5427_/B sky130_fd_sc_hd__nand2_1
X_5357_ _5357_/A _5357_/B vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__xnor2_2
XFILLER_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4308_ _4324_/C _4308_/B vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__xor2_1
X_5288_ _5486_/B vssd1 vssd1 vccd1 vccd1 _5485_/B sky130_fd_sc_hd__clkbuf_2
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4240_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6115__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5673__B _5675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6520__39 vssd1 vssd1 vccd1 vccd1 _6520__39/HI _6520_/A sky130_fd_sc_hd__conb_1
XFILLER_78_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_662 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _5109_/A vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__clkbuf_2
X_3610_ _4731_/B _4820_/B vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5583__B _5630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3541_ _4898_/A _3762_/B _3532_/A _3540_/Y vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__a31o_1
XFILLER_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _6379_/Q _6263_/C vssd1 vssd1 vccd1 vccd1 _6261_/B sky130_fd_sc_hd__and2_1
X_3472_ _3471_/A _3471_/B _3471_/C vssd1 vssd1 vccd1 vccd1 _3536_/B sky130_fd_sc_hd__a21o_1
X_5211_ _5211_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _5212_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6191_ _6352_/Q _6197_/B vssd1 vssd1 vccd1 vccd1 _6192_/A sky130_fd_sc_hd__and2_1
X_5142_ _5142_/A vssd1 vssd1 vccd1 vccd1 _5142_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3831__B _4051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5073_ _5062_/A _5061_/B _3950_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__a2bb2o_1
X_4024_ _4115_/A vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5975_ _5951_/A _5972_/X _5973_/Y _3380_/A vssd1 vssd1 vccd1 vccd1 _5976_/B sky130_fd_sc_hd__a31o_1
X_4926_ _4926_/A _4926_/B vssd1 vssd1 vccd1 vccd1 _5134_/B sky130_fd_sc_hd__xor2_4
X_4857_ _4857_/A _4865_/A vssd1 vssd1 vccd1 vccd1 _4857_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3808_ _3808_/A _3808_/B vssd1 vssd1 vccd1 vccd1 _3810_/C sky130_fd_sc_hd__xnor2_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6527_ _6527_/A _3236_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_4788_ _3494_/A _4787_/B _4787_/C _4787_/A vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__a22o_1
X_3739_ _3739_/A _3739_/B vssd1 vssd1 vccd1 vccd1 _3740_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3294__A _3294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5409_ _5409_/A _5409_/B vssd1 vssd1 vccd1 vccd1 _5535_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5768__C1 _6259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5859__A _5980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5760_ _5773_/A _5757_/Y _5759_/X _5815_/A vssd1 vssd1 vccd1 vccd1 _5760_/X sky130_fd_sc_hd__o22a_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _3661_/A _4675_/C _4785_/D _4645_/B vssd1 vssd1 vccd1 vccd1 _4712_/B sky130_fd_sc_hd__a22oi_1
X_5691_ _5691_/A _5935_/A _5691_/C _5691_/D vssd1 vssd1 vccd1 vccd1 _5819_/A sky130_fd_sc_hd__nor4_2
X_4642_ _4768_/D vssd1 vssd1 vccd1 vccd1 _4785_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_551 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4573_ _5001_/A vssd1 vssd1 vccd1 vccd1 _5714_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4003__A _4062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6312_ _6384_/CLK _6312_/D vssd1 vssd1 vccd1 vccd1 _6312_/Q sky130_fd_sc_hd__dfxtp_1
X_3524_ _3516_/Y _3529_/B _3526_/C vssd1 vssd1 vccd1 vccd1 _3525_/B sky130_fd_sc_hd__and3b_1
X_6243_ _6372_/Q _6239_/B _6242_/Y vssd1 vssd1 vccd1 vccd1 _6372_/D sky130_fd_sc_hd__o21a_1
X_3455_ _6298_/Q vssd1 vssd1 vccd1 vccd1 _6016_/A sky130_fd_sc_hd__clkbuf_2
X_6174_ _6346_/Q _6176_/B vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__and2_1
X_3386_ _3386_/A vssd1 vssd1 vccd1 vccd1 _3387_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5125_ _5125_/A _5125_/B _5125_/C vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__nand3_1
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5056_/A _5056_/B _5056_/C vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__or3_1
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4007_ _4007_/A _4007_/B _4007_/C vssd1 vssd1 vccd1 vccd1 _4008_/C sky130_fd_sc_hd__or3_1
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5958_ _5959_/A _5959_/C _5959_/B vssd1 vssd1 vccd1 vccd1 _5958_/Y sky130_fd_sc_hd__a21oi_1
X_4909_ _5203_/B _5203_/C _5203_/A vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__a21bo_1
X_5889_ _6098_/A vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__buf_2
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5009__A _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4583__A _4583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3199__A _3201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6383_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3258_/A vssd1 vssd1 vccd1 vccd1 _3245_/A sky130_fd_sc_hd__buf_6
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5812_ _6375_/Q _5776_/Y _5782_/X _5811_/X _6259_/A vssd1 vssd1 vccd1 vccd1 _6537_/A
+ sky130_fd_sc_hd__a221oi_2
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5743_ _5739_/X _5741_/Y _6214_/B vssd1 vssd1 vccd1 vccd1 _5743_/X sky130_fd_sc_hd__a21o_1
X_5674_ _5677_/A _5677_/B _5576_/Y _5581_/X vssd1 vssd1 vccd1 vccd1 _5674_/Y sky130_fd_sc_hd__o22ai_2
X_4625_ _5735_/B _5747_/A _5717_/A _5724_/A _5735_/A vssd1 vssd1 vccd1 vccd1 _5710_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4556_ _5698_/A _4563_/B _4555_/X vssd1 vssd1 vccd1 vccd1 _4556_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3507_ _3631_/A _3502_/X _3668_/A _3506_/X vssd1 vssd1 vccd1 vccd1 _3507_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5771__B _6061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4487_ _4487_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4488_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6226_ _6365_/Q _6227_/C _6225_/Y vssd1 vssd1 vccd1 vccd1 _6365_/D sky130_fd_sc_hd__o21a_1
X_3438_ _3549_/B vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_103_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3369_ _3690_/A vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__clkbuf_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6338_/Q _6337_/Q _6340_/Q _6339_/Q vssd1 vssd1 vccd1 vccd1 _6157_/X sky130_fd_sc_hd__and4_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5108_ _5108_/A _5104_/A vssd1 vssd1 vccd1 vccd1 _5109_/C sky130_fd_sc_hd__or2b_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6088_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__or2_1
X_5039_ _5001_/A _5183_/B _5038_/C vssd1 vssd1 vccd1 vccd1 _5040_/B sky130_fd_sc_hd__a21oi_1
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6562__78 vssd1 vssd1 vccd1 vccd1 _6562__78/HI _6562_/A sky130_fd_sc_hd__conb_1
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _6275_/Q _4410_/B vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5872__A _6187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5390_ _5390_/A _5390_/B vssd1 vssd1 vccd1 vccd1 _5401_/A sky130_fd_sc_hd__xnor2_1
XFILLER_98_112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4341_ _4341_/A _4341_/B vssd1 vssd1 vccd1 vccd1 _4374_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3392__A _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4272_ _4272_/A _4272_/B vssd1 vssd1 vccd1 vccd1 _4297_/A sky130_fd_sc_hd__xor2_2
X_3223_ _3226_/A vssd1 vssd1 vccd1 vccd1 _3223_/Y sky130_fd_sc_hd__inv_2
X_6011_ _6011_/A _6011_/B vssd1 vssd1 vccd1 vccd1 _6012_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4625__C1 _5724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3987_ _5097_/A _3987_/B vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5726_ _5737_/B _5737_/C _5737_/A vssd1 vssd1 vccd1 vccd1 _5792_/A sky130_fd_sc_hd__a21oi_1
X_5657_ _5885_/A _5657_/B vssd1 vssd1 vccd1 vccd1 _5657_/Y sky130_fd_sc_hd__xnor2_1
X_4608_ _4613_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4608_/X sky130_fd_sc_hd__and2_1
X_5588_ _5711_/A _5630_/A vssd1 vssd1 vccd1 vccd1 _5669_/B sky130_fd_sc_hd__xor2_1
X_4539_ _5724_/A _4583_/A vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6209_ _6360_/Q vssd1 vssd1 vccd1 vccd1 _6214_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5957__A _5957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5692__A _5819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5647__A1 _4138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3940__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3910_ _3922_/A _4484_/C vssd1 vssd1 vccd1 vccd1 _3923_/C sky130_fd_sc_hd__xor2_1
X_4890_ _4891_/A _4890_/B _4890_/C vssd1 vssd1 vccd1 vccd1 _4908_/A sky130_fd_sc_hd__nand3_1
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3841_ _4091_/B vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__clkbuf_2
X_3772_ _3772_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _3773_/B sky130_fd_sc_hd__and2_1
XFILLER_80_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6560_ _6560_/A _3320_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XANTENNA__3387__A _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5511_ _5865_/A _5511_/B _5512_/B vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__or3_1
X_6491_ _6491_/A _3192_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
X_6526__45 vssd1 vssd1 vccd1 vccd1 _6526__45/HI _6526_/A sky130_fd_sc_hd__conb_1
X_5442_ _5485_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5445_/B sky130_fd_sc_hd__and3_1
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5373_ _5373_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _5373_/X sky130_fd_sc_hd__or2b_1
XANTENNA__6210__B _6254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4324_ _5355_/A _4324_/B _4324_/C vssd1 vssd1 vccd1 vccd1 _4324_/Y sky130_fd_sc_hd__nand3_1
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5638__A1 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4255_ _4261_/A _4261_/B _4254_/X vssd1 vssd1 vccd1 vccd1 _4257_/B sky130_fd_sc_hd__a21boi_4
X_3206_ _3208_/A vssd1 vssd1 vccd1 vccd1 _3206_/Y sky130_fd_sc_hd__inv_2
X_4186_ _5320_/A _4268_/B vssd1 vssd1 vccd1 vccd1 _4187_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3297__A _3300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5709_ _5899_/A vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6595__TE_B _3319_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4856__A _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_30 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4591__A _4603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3654__B _3693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _4040_/A _4040_/B vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__xor2_1
XFILLER_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_516 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5991_ _5995_/A _5988_/X _5990_/Y vssd1 vssd1 vccd1 vccd1 _6294_/D sky130_fd_sc_hd__o21a_1
X_4942_ _4942_/A _4941_/Y vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__or2b_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4873_ _4873_/A _4873_/B _4873_/C vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__nand3_2
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3824_ _3734_/B _3764_/A _3764_/B _3823_/Y vssd1 vssd1 vccd1 vccd1 _3825_/B sky130_fd_sc_hd__o31ai_4
X_3755_ _5064_/A _3947_/B _3948_/B vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__and3_1
X_6543_ _6543_/A _3255_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_3686_ _3686_/A _3686_/B vssd1 vssd1 vccd1 vccd1 _3729_/A sky130_fd_sc_hd__nand2_1
X_5425_ _5425_/A _5425_/B vssd1 vssd1 vccd1 vccd1 _5449_/B sky130_fd_sc_hd__or2_1
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5356_ _4053_/A _5158_/B _5354_/A _5355_/X vssd1 vssd1 vccd1 vccd1 _5379_/A sky130_fd_sc_hd__a31o_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5287_ _5450_/B _5489_/B vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__nand2_1
X_4307_ _5426_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4238_ _4238_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__xnor2_2
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4169_ _4167_/Y _4168_/X _5404_/A _4207_/B vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__o211a_1
XFILLER_83_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6115__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3755__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4586__A _5646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_674 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6490__9 vssd1 vssd1 vccd1 vccd1 _6490__9/HI _6490_/A sky130_fd_sc_hd__conb_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3540_ _3540_/A _3540_/B vssd1 vssd1 vccd1 vccd1 _3540_/Y sky130_fd_sc_hd__nor2_1
X_5210_ _5211_/A _5211_/B vssd1 vssd1 vccd1 vccd1 _5212_/A sky130_fd_sc_hd__and2_1
X_3471_ _3471_/A _3471_/B _3471_/C vssd1 vssd1 vccd1 vccd1 _3536_/A sky130_fd_sc_hd__nand3_2
X_6190_ _6190_/A vssd1 vssd1 vccd1 vccd1 _6352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5141_ _5141_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__and3_1
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5072_ _5013_/A _5215_/B _5086_/B _5071_/A vssd1 vssd1 vccd1 vccd1 _5074_/B sky130_fd_sc_hd__a31o_1
XFILLER_69_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4023_ _5165_/A _4334_/B vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__nand2_2
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6216__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5974_ _3380_/A _5929_/A _5972_/X _5973_/Y _6244_/A vssd1 vssd1 vccd1 vccd1 _5974_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_100_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4925_ _4925_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4947_/A sky130_fd_sc_hd__nand2_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4856_ _4856_/A _4850_/B vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__or2b_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3807_ _4692_/A _3807_/B _3807_/C vssd1 vssd1 vccd1 vccd1 _3808_/B sky130_fd_sc_hd__and3_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6526_ _6526_/A _3235_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
XANTENNA__3575__A _3601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4787_ _4787_/A _4787_/B _4787_/C vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__and3_1
X_3738_ _3807_/C _3738_/B vssd1 vssd1 vccd1 vccd1 _3740_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3669_ _3668_/B _3668_/C _3668_/A vssd1 vssd1 vccd1 vccd1 _3672_/B sky130_fd_sc_hd__o21ai_1
XFILLER_69_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5408_ _5537_/B _5408_/B vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__xnor2_2
X_5339_ _5339_/A _5339_/B vssd1 vssd1 vccd1 vccd1 _5343_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5030__A _5196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_298 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5205__A _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6314__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3379__B _5957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4766_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _4719_/B sky130_fd_sc_hd__nand2_1
X_6568__84 vssd1 vssd1 vccd1 vccd1 _6568__84/HI _6568_/A sky130_fd_sc_hd__conb_1
XANTENNA__5875__A _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5690_ _5690_/A _5690_/B vssd1 vssd1 vccd1 vccd1 _5699_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _4768_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4572_ _5634_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4572_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4003__B _4051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6311_ _6357_/CLK _6311_/D vssd1 vssd1 vccd1 vccd1 _6311_/Q sky130_fd_sc_hd__dfxtp_1
X_3523_ _3522_/A _3522_/B _3529_/A _3522_/D vssd1 vssd1 vccd1 vccd1 _3526_/C sky130_fd_sc_hd__a22o_1
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6242_ _6242_/A _6248_/C vssd1 vssd1 vccd1 vccd1 _6242_/Y sky130_fd_sc_hd__nor2_1
X_3454_ _3522_/A vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173_ _6173_/A vssd1 vssd1 vccd1 vccd1 _6346_/D sky130_fd_sc_hd__clkbuf_1
X_3385_ _6304_/Q vssd1 vssd1 vccd1 vccd1 _3386_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _5388_/B vssd1 vssd1 vccd1 vccd1 _5158_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5055_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _5562_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _4018_/A _4006_/B vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__and2_1
XFILLER_72_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5769__B _6061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5957_ _5957_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__xor2_1
X_4908_ _4908_/A _4908_/B _4908_/C vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_530 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5888_ _5715_/A _5857_/X _5887_/Y _5872_/X vssd1 vssd1 vccd1 vccd1 _6277_/D sky130_fd_sc_hd__o211a_1
X_4839_ _4833_/A _4832_/C _4832_/B vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4725__A1 _4726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6509_ _6509_/A _3214_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5811_ _5806_/Y _5809_/X _5810_/X vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5742_ _6361_/Q vssd1 vssd1 vccd1 vccd1 _6214_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5673_ _5675_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5677_/B sky130_fd_sc_hd__xnor2_1
X_4624_ _4624_/A vssd1 vssd1 vccd1 vccd1 _5717_/A sky130_fd_sc_hd__inv_2
XFILLER_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4555_ _4555_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__and2_1
X_3506_ _3505_/A _3733_/A _3505_/C vssd1 vssd1 vccd1 vccd1 _3506_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5771__C _6061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4486_ _4486_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _4496_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5132__A1 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6225_ _6242_/A _6225_/B vssd1 vssd1 vccd1 vccd1 _6225_/Y sky130_fd_sc_hd__nor2_1
X_3437_ _3559_/B vssd1 vssd1 vccd1 vccd1 _3601_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3368_ _3520_/B vssd1 vssd1 vccd1 vccd1 _3690_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6156_/A vssd1 vssd1 vccd1 vccd1 _6340_/D sky130_fd_sc_hd__clkbuf_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5107_ _5107_/A _5107_/B _5107_/C vssd1 vssd1 vccd1 vccd1 _5113_/A sky130_fd_sc_hd__and3_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3299_/Y sky130_fd_sc_hd__inv_2
X_6087_ _6309_/Q _6310_/Q _6312_/Q _6311_/Q vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__or4_1
X_5038_ _5059_/A _5038_/B _5038_/C vssd1 vssd1 vccd1 vccd1 _5040_/A sky130_fd_sc_hd__and3_1
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4340_ _5484_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4341_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ _5358_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4272_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3222_ _3226_/A vssd1 vssd1 vccd1 vccd1 _3222_/Y sky130_fd_sc_hd__inv_2
X_6010_ _6003_/A _6003_/B _6001_/A vssd1 vssd1 vccd1 vccd1 _6011_/B sky130_fd_sc_hd__o21ai_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3986_ _5215_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5725_ _5671_/Y _5674_/Y _5749_/A _5677_/Y vssd1 vssd1 vccd1 vccd1 _5737_/C sky130_fd_sc_hd__o211ai_1
X_5656_ _5646_/Y _5651_/X _5655_/X vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__a21oi_1
X_4607_ _5605_/A _4548_/C _4548_/B vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__a21boi_1
X_5587_ _5679_/A _5637_/A vssd1 vssd1 vccd1 vccd1 _5669_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4538_ _4538_/A _4538_/B vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__xnor2_4
X_4469_ _4469_/A _4469_/B vssd1 vssd1 vccd1 vccd1 _4469_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6208_ _6354_/Q _6352_/D _6204_/X _6207_/X _5861_/X vssd1 vssd1 vccd1 vccd1 _6359_/D
+ sky130_fd_sc_hd__a32o_1
X_6139_ _5904_/X _6134_/X _6135_/X _6138_/X vssd1 vssd1 vccd1 vccd1 _6332_/D sky130_fd_sc_hd__a31o_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3419__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_411 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6586__102 vssd1 vssd1 vccd1 vccd1 _6586__102/HI _6586_/A sky130_fd_sc_hd__conb_1
XFILLER_96_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _3840_/A _3840_/B vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__xnor2_1
X_3771_ _3772_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5510_ _5510_/A _5510_/B vssd1 vssd1 vccd1 vccd1 _5512_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6490_ _6490_/A _3191_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
X_5441_ _5451_/A _5452_/B _5451_/B vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__o21ba_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5372_ _5373_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _5380_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4323_ _4323_/A _4323_/B vssd1 vssd1 vccd1 vccd1 _4323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _4254_/A _4253_/A vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__or2b_1
X_4185_ _4185_/A _4185_/B vssd1 vssd1 vccd1 vccd1 _4187_/A sky130_fd_sc_hd__xor2_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3205_ _3208_/A vssd1 vssd1 vccd1 vccd1 _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ _4492_/A _3969_/B vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__nand2_2
X_5708_ _6366_/Q _5707_/X _5697_/Y _6367_/Q vssd1 vssd1 vccd1 vccd1 _5708_/X sky130_fd_sc_hd__o22a_1
XFILLER_109_516 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4129__A2 _4168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5639_ _5639_/A _5639_/B vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__or2_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5033__A _5196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3812__A1 _5957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5990_ _5995_/A _6057_/A _5952_/X vssd1 vssd1 vccd1 vccd1 _5990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4941_ _4941_/A _4941_/B vssd1 vssd1 vccd1 vccd1 _4941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4872_ _4870_/A _4870_/B _4889_/A vssd1 vssd1 vccd1 vccd1 _4873_/C sky130_fd_sc_hd__a21o_1
X_3823_ _4933_/A _3503_/B _3764_/B _3822_/X vssd1 vssd1 vccd1 vccd1 _3823_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542_ _6542_/A _3254_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
X_3754_ _3754_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__xnor2_1
X_3685_ _3623_/A _3623_/B _3673_/B _3640_/X vssd1 vssd1 vccd1 vccd1 _3717_/C sky130_fd_sc_hd__a211o_1
XFILLER_106_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5424_ _5330_/A _5510_/B _5394_/B vssd1 vssd1 vccd1 vccd1 _5425_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5355_ _5355_/A _5355_/B _5359_/A vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__and3_1
X_5286_ _5286_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5297_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4306_ _4306_/A _4306_/B vssd1 vssd1 vccd1 vccd1 _4324_/C sky130_fd_sc_hd__xnor2_1
XFILLER_59_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4237_ _4237_/A _4237_/B vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3580__B _4898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4168_ _5199_/A _4168_/B _4168_/C vssd1 vssd1 vccd1 vccd1 _4168_/X sky130_fd_sc_hd__and3_1
XFILLER_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6369_/CLK sky130_fd_sc_hd__clkbuf_16
X_4099_ _4138_/A _4063_/B _4093_/B _4098_/X vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__a31o_1
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3755__B _3947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5698__A _5698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3470_ _3514_/A _3514_/B _3515_/B vssd1 vssd1 vccd1 vccd1 _3471_/C sky130_fd_sc_hd__nor3_1
XFILLER_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _5138_/A _5138_/B _5179_/A vssd1 vssd1 vccd1 vccd1 _5141_/C sky130_fd_sc_hd__a21bo_1
XFILLER_36_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5071_ _5071_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _5086_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4022_ _4022_/A _4071_/A vssd1 vssd1 vccd1 vccd1 _4334_/B sky130_fd_sc_hd__xor2_2
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_300 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5973_ _5691_/A _5967_/X _5949_/X vssd1 vssd1 vccd1 vccd1 _5973_/Y sky130_fd_sc_hd__o21ai_1
X_4924_ _5099_/A vssd1 vssd1 vccd1 vccd1 _5013_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4855_ _4855_/A _4855_/B _4855_/C vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__and3_1
X_3806_ _4698_/A _3502_/X _3734_/B _4933_/A vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__a22o_1
X_4786_ _4786_/A _4786_/B _4827_/A vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__nand3_1
X_6525_ _6525_/A _3232_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_3737_ _4796_/A _3700_/B _3697_/C _4645_/B vssd1 vssd1 vccd1 vccd1 _3738_/B sky130_fd_sc_hd__a22o_1
XFILLER_109_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3668_ _3668_/A _3668_/B _3668_/C vssd1 vssd1 vccd1 vccd1 _3672_/A sky130_fd_sc_hd__or3_1
X_5407_ _5403_/A _5403_/B _5406_/X vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__o21a_1
X_3599_ _3599_/A _3599_/B vssd1 vssd1 vccd1 vccd1 _3605_/B sky130_fd_sc_hd__xnor2_1
X_5338_ _5357_/A _5357_/B _5337_/X vssd1 vssd1 vccd1 vccd1 _5343_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5269_ _5269_/A vssd1 vssd1 vccd1 vccd1 _5444_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_480 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5205__B _5469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4640_ _4675_/C vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6583__99 vssd1 vssd1 vccd1 vccd1 _6583__99/HI _6583_/A sky130_fd_sc_hd__conb_1
X_4571_ _4569_/A _4569_/B _4570_/X vssd1 vssd1 vccd1 vccd1 _4571_/Y sky130_fd_sc_hd__a21oi_1
X_6310_ _6384_/CLK _6310_/D vssd1 vssd1 vccd1 vccd1 _6310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3522_ _3522_/A _3522_/B _3529_/A _3522_/D vssd1 vssd1 vccd1 vccd1 _3529_/B sky130_fd_sc_hd__nand4_1
X_6241_ _6372_/Q _6241_/B _6241_/C vssd1 vssd1 vccd1 vccd1 _6248_/C sky130_fd_sc_hd__and3_1
X_3453_ _3452_/A _3452_/B _3514_/A vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4300__A _6278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6172_ _6345_/Q _6176_/B vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__and2_1
X_5123_ _5123_/A _5123_/B vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__xor2_1
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3384_ _3384_/A vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5054_ _5554_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__and2_1
X_4005_ _4005_/A _4005_/B _4005_/C vssd1 vssd1 vccd1 vccd1 _4006_/B sky130_fd_sc_hd__or3_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6289__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4970__A _5145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _5943_/A _5943_/B _5691_/C _5957_/B vssd1 vssd1 vccd1 vccd1 _5959_/C sky130_fd_sc_hd__a2bb2o_1
X_4907_ _5247_/A _5290_/A vssd1 vssd1 vccd1 vccd1 _5203_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5887_ _5910_/A _5887_/B vssd1 vssd1 vccd1 vccd1 _5887_/Y sky130_fd_sc_hd__nand2_1
X_4838_ _4838_/A _4838_/B vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4725__A2 _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4769_ _4877_/B _4769_/B vssd1 vssd1 vccd1 vccd1 _4770_/C sky130_fd_sc_hd__nand2_1
X_6508_ _6508_/A _3213_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_96_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5913__A1 _5906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3943__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5810_ _6373_/Q _5808_/X _5781_/X _6374_/Q vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__a22o_1
XFILLER_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5741_ _5741_/A _5741_/B vssd1 vssd1 vccd1 vccd1 _5741_/Y sky130_fd_sc_hd__nand2_1
X_5672_ _5672_/A _5703_/A vssd1 vssd1 vccd1 vccd1 _5677_/A sky130_fd_sc_hd__or2b_1
XFILLER_30_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4623_ _5746_/B _5746_/C _5746_/A vssd1 vssd1 vccd1 vccd1 _5747_/A sky130_fd_sc_hd__a21o_1
X_4554_ _4555_/A _4555_/B vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__xor2_1
XFILLER_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3505_ _3505_/A _3733_/A _3505_/C vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__nand3_1
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4485_ _4486_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__and2_1
X_6224_ _6365_/Q _6227_/C vssd1 vssd1 vccd1 vccd1 _6225_/B sky130_fd_sc_hd__and2_1
XFILLER_103_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3436_ _3436_/A _3436_/B vssd1 vssd1 vccd1 vccd1 _3559_/B sky130_fd_sc_hd__and2_1
XFILLER_106_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6339_/Q _6165_/B vssd1 vssd1 vccd1 vccd1 _6156_/A sky130_fd_sc_hd__and2_1
X_3367_ _6289_/Q vssd1 vssd1 vccd1 vccd1 _3520_/B sky130_fd_sc_hd__clkbuf_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5106_ _5107_/A _5107_/B _5107_/C vssd1 vssd1 vccd1 vccd1 _5106_/Y sky130_fd_sc_hd__nand3_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6305_/Q _6306_/Q _6307_/Q _6308_/Q vssd1 vssd1 vccd1 vccd1 _6088_/A sky130_fd_sc_hd__or4_1
X_3298_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3298_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5037_/A _5059_/B vssd1 vssd1 vccd1 vccd1 _5038_/C sky130_fd_sc_hd__and2_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5939_ _3381_/B _5930_/X _5938_/Y _5872_/X vssd1 vssd1 vccd1 vccd1 _6285_/D sky130_fd_sc_hd__o211a_1
XANTENNA__6304__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6139__A1 _5904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6553__69 vssd1 vssd1 vccd1 vccd1 _6553__69/HI _6553_/A sky130_fd_sc_hd__conb_1
XANTENNA__4769__B _4769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A _4270_/B vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__or2_1
X_3221_ _3227_/A vssd1 vssd1 vccd1 vccd1 _3226_/A sky130_fd_sc_hd__buf_6
XFILLER_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3985_ _5199_/A vssd1 vssd1 vccd1 vccd1 _5215_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5724_ _5724_/A _5793_/A vssd1 vssd1 vccd1 vccd1 _5724_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_10_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5655_ _5653_/Y _5651_/C _5651_/B _5654_/Y vssd1 vssd1 vccd1 vccd1 _5655_/X sky130_fd_sc_hd__o211a_1
X_4606_ _4621_/B _4606_/B vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__xnor2_1
X_5586_ _5586_/A _5586_/B vssd1 vssd1 vccd1 vccd1 _5637_/A sky130_fd_sc_hd__xnor2_4
X_4537_ _4537_/A _4537_/B vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__xor2_4
X_4468_ _4523_/A _4523_/B _4467_/Y vssd1 vssd1 vccd1 vccd1 _4518_/B sky130_fd_sc_hd__a21o_2
X_6207_ _6353_/Q _6205_/X _6206_/X _6359_/Q vssd1 vssd1 vccd1 vccd1 _6207_/X sky130_fd_sc_hd__o31a_1
X_3419_ _3387_/A _3391_/A _6300_/Q vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__a21o_2
X_4399_ _4399_/A _4399_/B vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__xor2_1
X_6138_ _6325_/Q _6324_/Q _6137_/X _6282_/D vssd1 vssd1 vccd1 vccd1 _6138_/X sky130_fd_sc_hd__o31a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6069_ _6306_/Q _6073_/B vssd1 vssd1 vccd1 vccd1 _6070_/A sky130_fd_sc_hd__and2_1
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5041__B2 _5145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4607__A1 _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_607 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3770_ _3735_/A _3774_/A _3741_/B _3740_/B _3740_/A vssd1 vssd1 vccd1 vccd1 _3772_/B
+ sky130_fd_sc_hd__a32oi_1
XFILLER_9_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5440_ _5440_/A _5440_/B _5440_/C vssd1 vssd1 vccd1 vccd1 _5451_/B sky130_fd_sc_hd__and3_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6060__A _6060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5371_ _5390_/A _5390_/B _5370_/X vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__a21bo_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _4322_/A _4322_/B vssd1 vssd1 vccd1 vccd1 _4329_/B sky130_fd_sc_hd__xnor2_2
X_4253_ _4253_/A _4254_/A vssd1 vssd1 vccd1 vccd1 _4261_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5404__A _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3204_ _3208_/A vssd1 vssd1 vccd1 vccd1 _3204_/Y sky130_fd_sc_hd__inv_2
X_4184_ _5231_/A _4367_/B vssd1 vssd1 vccd1 vccd1 _4185_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6384_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4962__B _5013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_412 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3968_ _4479_/B _3968_/B vssd1 vssd1 vccd1 vccd1 _3969_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5906_/A _5700_/X _5705_/X _5706_/X vssd1 vssd1 vccd1 vccd1 _5707_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6517__36 vssd1 vssd1 vccd1 vccd1 _6517__36/HI _6517_/A sky130_fd_sc_hd__conb_1
X_3899_ _3938_/A _3938_/B _3938_/C vssd1 vssd1 vccd1 vccd1 _4479_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5638_ _5714_/A _5657_/B _5637_/Y vssd1 vssd1 vccd1 vccd1 _5639_/B sky130_fd_sc_hd__a21oi_1
X_5569_ _5559_/A _5559_/B _5568_/X vssd1 vssd1 vccd1 vccd1 _5675_/A sky130_fd_sc_hd__a21oi_4
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5314__A _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6211__B1 _5952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_550 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6531__50 vssd1 vssd1 vccd1 vccd1 _6531__50/HI _6531_/A sky130_fd_sc_hd__conb_1
XFILLER_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4940_ _4941_/A _4941_/B vssd1 vssd1 vccd1 vccd1 _4942_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4871_ _4865_/A _4885_/A _4867_/A _4867_/B vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__o22ai_2
X_3822_ _3380_/A _3502_/X _3503_/A vssd1 vssd1 vccd1 vccd1 _3822_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6541_ _6541_/A _3253_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
X_3753_ _5011_/A _4168_/B vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__nand2_1
X_3684_ _3672_/A _3672_/B _3672_/C vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__a21o_1
X_5423_ _5484_/C vssd1 vssd1 vccd1 vccd1 _5510_/B sky130_fd_sc_hd__clkbuf_2
X_5354_ _5354_/A _5354_/B vssd1 vssd1 vccd1 vccd1 _5359_/A sky130_fd_sc_hd__xnor2_1
XFILLER_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _4334_/A _4337_/B _4337_/C vssd1 vssd1 vccd1 vccd1 _4306_/B sky130_fd_sc_hd__and3_1
X_5285_ _5285_/A _5285_/B vssd1 vssd1 vccd1 vccd1 _5318_/A sky130_fd_sc_hd__xnor2_2
X_4236_ _4236_/A _4236_/B vssd1 vssd1 vccd1 vccd1 _4261_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4167_ _4167_/A _4167_/B vssd1 vssd1 vccd1 vccd1 _4167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ _5109_/A _4138_/B _4098_/C vssd1 vssd1 vccd1 vccd1 _4098_/X sky130_fd_sc_hd__and3_1
XFILLER_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5070_ _5070_/A _5070_/B vssd1 vssd1 vccd1 vccd1 _5071_/B sky130_fd_sc_hd__and2_1
X_4021_ _4021_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4031_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5972_ _5691_/A _3379_/A _5959_/X _5966_/B vssd1 vssd1 vccd1 vccd1 _5972_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3202__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4923_ _4923_/A _4923_/B vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__xor2_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4854_ _4854_/A _4870_/A vssd1 vssd1 vccd1 vccd1 _4855_/C sky130_fd_sc_hd__nand2_1
X_3805_ _3805_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _3810_/A sky130_fd_sc_hd__or2_1
X_4785_ _4785_/A _4846_/A _4785_/C _4785_/D vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__nand4_1
XANTENNA__6232__B _6254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3736_ _3763_/A _3762_/B vssd1 vssd1 vccd1 vccd1 _3807_/C sky130_fd_sc_hd__nand2_1
X_6524_ _6524_/A _3231_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_109_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3667_ _3686_/B _3665_/X _3508_/A _3508_/Y vssd1 vssd1 vccd1 vccd1 _3668_/C sky130_fd_sc_hd__a211oi_1
X_5406_ _5409_/B _5409_/A vssd1 vssd1 vccd1 vccd1 _5406_/X sky130_fd_sc_hd__or2b_1
X_3598_ _3592_/X _3598_/B vssd1 vssd1 vccd1 vccd1 _3599_/B sky130_fd_sc_hd__and2b_1
X_5337_ _5336_/B _5337_/B vssd1 vssd1 vccd1 vccd1 _5337_/X sky130_fd_sc_hd__and2b_1
XFILLER_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5268_ _5268_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5544_/B sky130_fd_sc_hd__xnor2_2
X_4219_ _4213_/A _4212_/B _4212_/A vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__o21ba_2
X_5199_ _5199_/A _5316_/B vssd1 vssd1 vccd1 vccd1 _5200_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4976__B1 _4961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6501__20 vssd1 vssd1 vccd1 vccd1 _6501__20/HI _6501_/A sky130_fd_sc_hd__conb_1
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4431__A2 _4153_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4570_ _5899_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4570_/X sky130_fd_sc_hd__and2_1
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ _6288_/Q _3436_/A _3436_/B _3556_/B _6289_/Q vssd1 vssd1 vccd1 vccd1 _3522_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6240_ _6241_/B _6241_/C _6239_/Y vssd1 vssd1 vccd1 vccd1 _6371_/D sky130_fd_sc_hd__o21a_1
X_3452_ _3452_/A _3452_/B _3514_/A vssd1 vssd1 vccd1 vccd1 _3465_/A sky130_fd_sc_hd__nand3_1
XFILLER_115_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6171_ _6171_/A vssd1 vssd1 vccd1 vccd1 _6345_/D sky130_fd_sc_hd__clkbuf_1
X_3383_ _3383_/A vssd1 vssd1 vccd1 vccd1 _3384_/A sky130_fd_sc_hd__clkbuf_2
X_5122_ _5104_/A _5104_/B _5104_/C vssd1 vssd1 vccd1 vccd1 _5141_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5554_/A _5054_/B vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4004_ _4005_/A _4005_/B _4005_/C vssd1 vssd1 vccd1 vccd1 _4018_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_646 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5955_ _5955_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__or2_1
X_6559__75 vssd1 vssd1 vccd1 vccd1 _6559__75/HI _6559_/A sky130_fd_sc_hd__conb_1
XFILLER_80_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4906_ _5289_/A _5289_/B vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__and2_1
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5886_ _5886_/A _5886_/B vssd1 vssd1 vccd1 vccd1 _5887_/B sky130_fd_sc_hd__xnor2_1
X_4837_ _4916_/B _4837_/B vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__xnor2_4
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4768_ _4842_/B _4864_/B _4768_/C _4768_/D vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__nand4_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4699_ _4937_/B _4699_/B vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__or2_1
X_6507_ _6507_/A _3212_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_3719_ _3718_/A _3718_/B _3718_/C _3718_/D vssd1 vssd1 vccd1 vccd1 _3720_/B sky130_fd_sc_hd__a22o_1
XANTENNA__4698__A _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6369_ _6369_/CLK _6369_/D vssd1 vssd1 vccd1 vccd1 _6369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_532 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _5741_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5576_/Y _5581_/X _5668_/X _5670_/X vssd1 vssd1 vccd1 vccd1 _5671_/Y sky130_fd_sc_hd__a22oi_2
X_4622_ _5735_/B _4622_/B vssd1 vssd1 vccd1 vccd1 _5746_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4553_ _4553_/A _4559_/A vssd1 vssd1 vccd1 vccd1 _4555_/B sky130_fd_sc_hd__xor2_1
X_4484_ _4548_/A _4484_/B _4484_/C vssd1 vssd1 vccd1 vccd1 _4486_/B sky130_fd_sc_hd__and3_1
X_3504_ _3464_/A _3464_/B _3463_/A vssd1 vssd1 vccd1 vccd1 _3505_/C sky130_fd_sc_hd__o21bai_2
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6223_ _6364_/Q _6218_/B _6222_/Y vssd1 vssd1 vccd1 vccd1 _6364_/D sky130_fd_sc_hd__o21a_1
X_3435_ _6290_/Q vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3366_ _4312_/A vssd1 vssd1 vccd1 vccd1 _5936_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6154_ _6154_/A vssd1 vssd1 vccd1 vccd1 _6339_/D sky130_fd_sc_hd__clkbuf_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5105_ _5103_/A _5103_/B _5141_/A vssd1 vssd1 vccd1 vccd1 _5107_/C sky130_fd_sc_hd__a21bo_1
X_3297_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3297_/Y sky130_fd_sc_hd__inv_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6492__11 vssd1 vssd1 vccd1 vccd1 _6492__11/HI _6492_/A sky130_fd_sc_hd__conb_1
X_6085_ _6305_/Q _6306_/Q _6307_/Q _6308_/Q vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__and4_1
X_5036_ _3903_/A _5180_/D _5065_/B _5035_/A vssd1 vssd1 vccd1 vccd1 _5042_/B sky130_fd_sc_hd__a31o_1
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5840__B2 _5733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5938_ _5936_/X _5937_/Y _5970_/A vssd1 vssd1 vccd1 vccd1 _5938_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5869_ _5866_/X _5867_/Y _5910_/A vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5831__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__B2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3300__A _3300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4115__B _4367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4131__A _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3220_ _3220_/A vssd1 vssd1 vccd1 vccd1 _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6359_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5897__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3984_ _3984_/A _3984_/B vssd1 vssd1 vccd1 vccd1 _4040_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3210__A _3214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4025__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5723_ _5735_/B _5747_/A _5735_/A vssd1 vssd1 vccd1 vccd1 _5793_/A sky130_fd_sc_hd__a21oi_2
XFILLER_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5654_ _5740_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5654_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3864__B _4138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4605_ _4605_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4611_/C sky130_fd_sc_hd__and2_1
X_5585_ _5585_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__xnor2_2
XFILLER_116_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4536_ _4536_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _4537_/B sky130_fd_sc_hd__nand2_1
X_4467_ _4467_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _4467_/Y sky130_fd_sc_hd__nor2_1
X_4398_ _4399_/A _4399_/B _4397_/X vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__o21ai_1
X_6206_ _6356_/Q _6355_/Q _6358_/Q _6357_/Q vssd1 vssd1 vccd1 vccd1 _6206_/X sky130_fd_sc_hd__or4_1
X_3418_ _6299_/Q _6298_/Q _3449_/A _4749_/A vssd1 vssd1 vccd1 vccd1 _3458_/A sky130_fd_sc_hd__or4_2
X_3349_ _4645_/B vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__buf_2
X_6137_ _6327_/Q _6326_/Q _6137_/C vssd1 vssd1 vccd1 vccd1 _6137_/X sky130_fd_sc_hd__or3_1
XANTENNA_input8_A la1_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6068_ _6068_/A vssd1 vssd1 vccd1 vccd1 _6306_/D sky130_fd_sc_hd__clkbuf_1
X_5019_ _5019_/A _5019_/B vssd1 vssd1 vccd1 vccd1 _5020_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5370_ _5370_/A _5370_/B _5369_/B vssd1 vssd1 vccd1 vccd1 _5370_/X sky130_fd_sc_hd__or3b_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4321_ _4350_/A _4350_/B _4320_/X vssd1 vssd1 vccd1 vccd1 _4322_/B sky130_fd_sc_hd__o21a_1
X_4252_ _4273_/A _4273_/B _4251_/A vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__o21a_1
X_3203_ _3227_/A vssd1 vssd1 vccd1 vccd1 _3208_/A sky130_fd_sc_hd__buf_8
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4183_ _5231_/B _4337_/B _4337_/C vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__and3_1
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3205__A _3208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6048__A1 _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4231__B1 _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3967_ _4479_/B _4479_/C _4479_/A vssd1 vssd1 vccd1 vccd1 _4521_/A sky130_fd_sc_hd__a21oi_1
X_5706_ _5841_/B vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3898_ _3919_/B _3898_/B vssd1 vssd1 vccd1 vccd1 _3938_/C sky130_fd_sc_hd__nand2_1
X_5637_ _5637_/A _5637_/B vssd1 vssd1 vccd1 vccd1 _5637_/Y sky130_fd_sc_hd__nor2_1
X_5568_ _5023_/B _5024_/A _4997_/B _5567_/Y vssd1 vssd1 vccd1 vccd1 _5568_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4519_ _5710_/A _4569_/A vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__or2b_1
X_5499_ _5499_/A _5527_/A vssd1 vssd1 vccd1 vccd1 _5529_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5314__B _5358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3785__A _3840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_562 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6317__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4870_ _4870_/A _4870_/B _4889_/A vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__nand3_2
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3821_ _3813_/A _3813_/B _3811_/A vssd1 vssd1 vccd1 vccd1 _3825_/A sky130_fd_sc_hd__a21o_2
XANTENNA__5005__A2 _4961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6540_ _6540_/A _3251_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _4207_/B vssd1 vssd1 vccd1 vccd1 _3947_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3683_ _5091_/A vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__xnor2_1
X_5353_ _5386_/A _5388_/B vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__nand2_1
X_4304_ _4317_/A _4317_/B _4303_/Y vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__a21oi_2
XFILLER_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ _5284_/A _5284_/B vssd1 vssd1 vccd1 vccd1 _5285_/A sky130_fd_sc_hd__or2_1
XFILLER_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4235_ _5278_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _4236_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5134__B _5134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4166_ _5355_/A _4166_/B vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__nand2_1
X_4097_ _4097_/A _4097_/B vssd1 vssd1 vccd1 vccd1 _4100_/B sky130_fd_sc_hd__xor2_1
XFILLER_82_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4999_ _5023_/B _4999_/B vssd1 vssd1 vccd1 vccd1 _5052_/A sky130_fd_sc_hd__or2_1
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5325__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4020_ _5158_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__nand2_1
XFILLER_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5971_ _5691_/A _5930_/X _5970_/Y _5945_/X vssd1 vssd1 vccd1 vccd1 _6290_/D sky130_fd_sc_hd__o211a_1
X_4922_ _4926_/A _4926_/B _4746_/A vssd1 vssd1 vccd1 vccd1 _4923_/B sky130_fd_sc_hd__a21o_2
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4853_ _4854_/A _4853_/B _4853_/C vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__nand3_1
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3804_ _3804_/A _3804_/B vssd1 vssd1 vccd1 vccd1 _3815_/A sky130_fd_sc_hd__nand2_1
X_4784_ _4771_/A _4770_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _4786_/B sky130_fd_sc_hd__a21o_1
X_6523_ _6523_/A _3230_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
X_3735_ _3735_/A _3774_/A vssd1 vssd1 vccd1 vccd1 _3741_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5405_ _5355_/A _5158_/B _5389_/A _5404_/X vssd1 vssd1 vccd1 vccd1 _5409_/A sky130_fd_sc_hd__a31o_1
X_3666_ _3508_/A _3508_/Y _3686_/B _3665_/X vssd1 vssd1 vccd1 vccd1 _3668_/B sky130_fd_sc_hd__o211a_1
X_3597_ _3617_/A _3617_/B _3617_/C vssd1 vssd1 vccd1 vccd1 _3627_/B sky130_fd_sc_hd__a21o_1
X_5336_ _5337_/B _5336_/B vssd1 vssd1 vccd1 vccd1 _5357_/B sky130_fd_sc_hd__xnor2_2
X_5267_ _5267_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5268_/B sky130_fd_sc_hd__xnor2_1
X_4218_ _4220_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__or2b_1
XFILLER_102_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5198_ _5198_/A _5198_/B vssd1 vssd1 vccd1 vccd1 _5215_/C sky130_fd_sc_hd__nor2_1
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5217__A2 _5013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4149_ _3614_/Y _4148_/X _3635_/B vssd1 vssd1 vccd1 vccd1 _4301_/B sky130_fd_sc_hd__o21ba_1
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4728__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3303__A _3306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3520_ _5995_/A _3520_/B _6288_/Q _5325_/B vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__nand4_1
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3451_ _6290_/Q _3477_/D _3522_/B vssd1 vssd1 vccd1 vccd1 _3514_/A sky130_fd_sc_hd__and3_1
XFILLER_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6170_ _6344_/Q _6176_/B vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__and2_1
X_3382_ _5715_/B vssd1 vssd1 vccd1 vccd1 _3383_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _5119_/A _5118_/C _5118_/A vssd1 vssd1 vccd1 vccd1 _5550_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5052_ _5052_/A _5052_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__xnor2_1
X_4003_ _4062_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4005_/C sky130_fd_sc_hd__and2_1
XFILLER_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3213__A _3214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5954_ _5955_/A _5951_/X _5953_/Y vssd1 vssd1 vccd1 vccd1 _6287_/D sky130_fd_sc_hd__o21a_1
X_4905_ _4905_/A _4905_/B vssd1 vssd1 vccd1 vccd1 _5289_/B sky130_fd_sc_hd__xnor2_1
X_5885_ _5885_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5886_/B sky130_fd_sc_hd__xnor2_1
X_4836_ _4838_/A _4838_/B _4835_/Y vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__o21a_1
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4767_ _4879_/B _4768_/C _4768_/D _4879_/A vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__a22o_1
X_6506_ _6506_/A _3211_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
X_4698_ _4698_/A _4931_/A _4698_/C vssd1 vssd1 vccd1 vccd1 _4699_/B sky130_fd_sc_hd__and3_1
X_3718_ _3718_/A _3718_/B _3718_/C _3718_/D vssd1 vssd1 vccd1 vccd1 _3782_/A sky130_fd_sc_hd__nand4_4
XFILLER_4_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3649_ _3649_/A _3649_/B _3649_/C vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__nand3_1
X_6368_ _6369_/CLK _6368_/D vssd1 vssd1 vccd1 vccd1 _6368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5319_ _5271_/X _5312_/X _5311_/X vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__a21bo_1
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6299_ _6345_/CLK _6299_/D vssd1 vssd1 vccd1 vccd1 _6299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6335_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3687__B _3693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5583_/X _5669_/Y _5584_/Y vssd1 vssd1 vccd1 vccd1 _5670_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4621_ _4621_/A _4621_/B vssd1 vssd1 vccd1 vccd1 _4622_/B sky130_fd_sc_hd__or2_1
XFILLER_30_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4799__A _4818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4552_ _5619_/A vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__buf_2
XFILLER_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4483_ _3937_/X _4492_/B _4491_/A vssd1 vssd1 vccd1 vccd1 _4490_/A sky130_fd_sc_hd__a21o_1
X_3503_ _3503_/A _3503_/B vssd1 vssd1 vccd1 vccd1 _3733_/A sky130_fd_sc_hd__and2_1
XANTENNA__3208__A _3208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3434_ _5935_/A _3432_/A _3807_/B _3474_/A vssd1 vssd1 vccd1 vccd1 _3513_/A sky130_fd_sc_hd__a31o_1
X_6222_ _6242_/A _6227_/C vssd1 vssd1 vccd1 vccd1 _6222_/Y sky130_fd_sc_hd__nor2_1
X_3365_ _3631_/A vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__clkbuf_1
X_6153_ _6338_/Q _6165_/B vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__and2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5104_/A _5104_/B _5104_/C vssd1 vssd1 vccd1 vccd1 _5141_/A sky130_fd_sc_hd__nand3_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3296_/Y sky130_fd_sc_hd__inv_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6309_/Q _6310_/Q _6312_/Q _6311_/Q vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__and4_1
X_5035_ _5035_/A _5035_/B vssd1 vssd1 vccd1 vccd1 _5065_/B sky130_fd_sc_hd__nor2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5937_ _5937_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5937_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3603__B2 _4882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5868_ _5868_/A vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4819_ _4822_/A _4819_/B vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__or2_1
X_5799_ _6369_/Q vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_468 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3983_ _3984_/A _3984_/B vssd1 vssd1 vccd1 vccd1 _4007_/A sky130_fd_sc_hd__and2_1
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ _5838_/B _5744_/C vssd1 vssd1 vccd1 vccd1 _5732_/A sky130_fd_sc_hd__nor2_1
X_5653_ _5740_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _5653_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4604_ _4605_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4611_/B sky130_fd_sc_hd__nor2_1
X_5584_ _5683_/A _5624_/A vssd1 vssd1 vccd1 vccd1 _5584_/Y sky130_fd_sc_hd__xnor2_1
X_4535_ _5735_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__or2b_1
XFILLER_7_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4466_ _4538_/A _4538_/B _4465_/X vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__a21o_2
XFILLER_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4397_ _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__or2_1
X_6205_ _6352_/Q _6351_/Q _6354_/Q vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__or3_1
X_3417_ _3469_/A _3469_/B _3416_/X vssd1 vssd1 vccd1 vccd1 _3432_/A sky130_fd_sc_hd__a21o_1
X_3348_ _3645_/B vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_503 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6136_ _6329_/Q _6328_/Q _6331_/Q _6330_/Q vssd1 vssd1 vccd1 vccd1 _6137_/C sky130_fd_sc_hd__or4_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_666 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6067_ _6305_/Q _6073_/B vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__and2_1
X_3279_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3279_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5018_ _5019_/A _5019_/B vssd1 vssd1 vccd1 vccd1 _5020_/A sky130_fd_sc_hd__or2_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5998__A _6000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3311__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6593__109 vssd1 vssd1 vccd1 vccd1 _6593__109/HI _6593_/A sky130_fd_sc_hd__conb_1
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4320_ _4320_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__or2b_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4251_ _4251_/A _4251_/B vssd1 vssd1 vccd1 vccd1 _4273_/B sky130_fd_sc_hd__nand2_1
X_3202_ input1/X vssd1 vssd1 vccd1 vccd1 _3227_/A sky130_fd_sc_hd__buf_2
XFILLER_101_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4182_ _4182_/A _4182_/B vssd1 vssd1 vccd1 vccd1 _4214_/B sky130_fd_sc_hd__xnor2_4
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3806__A1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3806__B2 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3966_ _4014_/A _4014_/B vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__and2_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5705_ _5773_/A _5702_/Y _5703_/Y _5815_/A vssd1 vssd1 vccd1 vccd1 _5705_/X sky130_fd_sc_hd__o22a_1
X_3897_ _3897_/A _3897_/B vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__nand2_1
X_5636_ _5637_/A _5637_/B vssd1 vssd1 vccd1 vccd1 _5657_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5567_ _4996_/A _4993_/Y _4995_/S vssd1 vssd1 vccd1 vccd1 _5567_/Y sky130_fd_sc_hd__a21oi_1
X_4518_ _4518_/A _4518_/B vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__xor2_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5498_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5527_/A sky130_fd_sc_hd__and2_1
X_4449_ _5514_/A _4449_/B vssd1 vssd1 vccd1 vccd1 _4581_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6119_ _6324_/Q _6127_/B vssd1 vssd1 vccd1 vccd1 _6120_/A sky130_fd_sc_hd__and2_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5330__B _5485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3785__B _3785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6508__27 vssd1 vssd1 vccd1 vccd1 _6508__27/HI _6508_/A sky130_fd_sc_hd__conb_1
XFILLER_6_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5505__B _5505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3306__A _3306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5789__B2 _5733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3820_ _3816_/B _3818_/B _3816_/A vssd1 vssd1 vccd1 vccd1 _3829_/B sky130_fd_sc_hd__a21bo_1
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _3987_/B vssd1 vssd1 vccd1 vccd1 _4207_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5961__A1 _5957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3682_ _5130_/A vssd1 vssd1 vccd1 vccd1 _5091_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5421_ _5421_/A _5421_/B vssd1 vssd1 vccd1 vccd1 _5429_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_3_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6522__41 vssd1 vssd1 vccd1 vccd1 _6522__41/HI _6522_/A sky130_fd_sc_hd__conb_1
X_5352_ _5348_/X _5362_/B _5361_/A vssd1 vssd1 vccd1 vccd1 _5354_/A sky130_fd_sc_hd__a21o_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4303_ _4303_/A _4332_/A vssd1 vssd1 vccd1 vccd1 _4303_/Y sky130_fd_sc_hd__nor2_1
X_5283_ _5301_/A _5301_/B vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__and2_1
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3216__A _3220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4234_ _4231_/X _4234_/B vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _4216_/B _4216_/A vssd1 vssd1 vccd1 vccd1 _4165_/X sky130_fd_sc_hd__and2b_1
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4106_/A _4106_/B _4095_/X vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__o21ai_1
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4998_ _4998_/A _4998_/B _4998_/C vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__nor3_1
XFILLER_11_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3949_ _3957_/A _3949_/B vssd1 vssd1 vccd1 vccd1 _3991_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5619_ _5619_/A _5619_/B vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5325__B _5325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5970_ _5970_/A _5970_/B vssd1 vssd1 vccd1 vccd1 _5970_/Y sky130_fd_sc_hd__nand2_1
X_4921_ _5008_/A _5008_/B _4920_/Y vssd1 vssd1 vccd1 vccd1 _4926_/B sky130_fd_sc_hd__a21o_1
X_4852_ _4869_/A _4852_/B _4852_/C vssd1 vssd1 vccd1 vccd1 _4853_/C sky130_fd_sc_hd__nand3b_1
X_3803_ _3950_/A vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4783_ _4783_/A _4783_/B vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6522_ _6522_/A _3321_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
X_3734_ _4634_/A _3734_/B _3734_/C vssd1 vssd1 vccd1 vccd1 _3774_/A sky130_fd_sc_hd__nand3_1
X_6499__18 vssd1 vssd1 vccd1 vccd1 _6499__18/HI _6499_/A sky130_fd_sc_hd__conb_1
X_3665_ _3686_/A _3664_/B _3664_/C vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5404_ _5404_/A _5404_/B _5404_/C vssd1 vssd1 vccd1 vccd1 _5404_/X sky130_fd_sc_hd__and3_1
XANTENNA__5145__B _5145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6384_ _6384_/CLK _6384_/D vssd1 vssd1 vccd1 vccd1 _6384_/Q sky130_fd_sc_hd__dfxtp_1
X_3596_ _3615_/B _3615_/A vssd1 vssd1 vccd1 vccd1 _3617_/C sky130_fd_sc_hd__and2b_1
X_5335_ _5360_/A _5360_/B _5334_/A vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__o21ba_1
XFILLER_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5266_ _5578_/A _5578_/B _5578_/C vssd1 vssd1 vccd1 vccd1 _5579_/A sky130_fd_sc_hd__o21ai_1
X_4217_ _4217_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__xnor2_1
X_5197_ _5195_/A _5358_/B _5158_/B _5133_/A vssd1 vssd1 vccd1 vccd1 _5198_/B sky130_fd_sc_hd__a22oi_1
XFILLER_56_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4148_ _3634_/B _3614_/B _3633_/X vssd1 vssd1 vccd1 vccd1 _4148_/X sky130_fd_sc_hd__a21bo_1
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4079_ _4079_/A _4207_/B vssd1 vssd1 vccd1 vccd1 _4082_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4505__A _4516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6307__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4728__A2 _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6357_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4416__A1 _4266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5246__A _5246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5144__A2 _5038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3450_ _3492_/A vssd1 vssd1 vccd1 vccd1 _3522_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3381_ _5691_/A _3381_/B _5691_/C _5691_/D vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__or4_4
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5120_ _5552_/B _5120_/B vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__xnor2_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5051_ _5056_/B _5056_/C _5056_/A vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__o21ai_1
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4053_/A vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5953_ _5955_/A _5951_/X _5952_/X vssd1 vssd1 vccd1 vccd1 _5953_/Y sky130_fd_sc_hd__a21oi_1
X_4904_ _4898_/A _4898_/B _3611_/A _4726_/A vssd1 vssd1 vccd1 vccd1 _4905_/B sky130_fd_sc_hd__o22a_1
X_5884_ _5899_/B vssd1 vssd1 vccd1 vccd1 _5906_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4835_ _4835_/A _4835_/B vssd1 vssd1 vccd1 vccd1 _4835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5907__A1 _5755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4766_ _4766_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__xnor2_1
X_3717_ _3717_/A _3717_/B _3717_/C vssd1 vssd1 vccd1 vccd1 _3718_/D sky130_fd_sc_hd__nand3_1
X_6505_ _6505_/A _3210_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_107_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4697_ _4698_/A _4931_/A _4698_/C vssd1 vssd1 vccd1 vccd1 _4937_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5135__A2 _5134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3648_ _3647_/B _3647_/C _3647_/A vssd1 vssd1 vccd1 vccd1 _3649_/C sky130_fd_sc_hd__o21ai_1
X_6367_ _6383_/CLK _6367_/D vssd1 vssd1 vccd1 vccd1 _6367_/Q sky130_fd_sc_hd__dfxtp_1
X_3579_ _4842_/A _4877_/D vssd1 vssd1 vccd1 vccd1 _4898_/B sky130_fd_sc_hd__nand2_2
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5318_ _5318_/A _5318_/B vssd1 vssd1 vccd1 vccd1 _5337_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6298_ _6335_/CLK _6298_/D vssd1 vssd1 vccd1 vccd1 _6298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5249_ _5328_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__and2_1
XFILLER_29_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4235__A _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3314__A _3318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4637__B2 _4814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4528_/X _4616_/X _4617_/X _4618_/Y _4619_/X vssd1 vssd1 vccd1 vccd1 _5746_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4551_ _4961_/A vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__buf_2
X_6564__80 vssd1 vssd1 vccd1 vccd1 _6564__80/HI _6564_/A sky130_fd_sc_hd__conb_1
X_4482_ _4482_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__nor2_1
X_3502_ _3697_/C vssd1 vssd1 vccd1 vccd1 _3502_/X sky130_fd_sc_hd__clkbuf_2
X_3433_ _3473_/A _3473_/B vssd1 vssd1 vccd1 vccd1 _3474_/A sky130_fd_sc_hd__and2_1
X_6221_ _6364_/Q _6363_/Q _6221_/C vssd1 vssd1 vccd1 vccd1 _6227_/C sky130_fd_sc_hd__and3_1
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6152_ _6152_/A vssd1 vssd1 vccd1 vccd1 _6338_/D sky130_fd_sc_hd__clkbuf_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5103_ _5103_/A _5103_/B vssd1 vssd1 vccd1 vccd1 _5104_/C sky130_fd_sc_hd__xor2_1
X_3364_ _4846_/A vssd1 vssd1 vccd1 vccd1 _3631_/A sky130_fd_sc_hd__clkbuf_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__buf_8
XANTENNA__3224__A _3226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6083_/A vssd1 vssd1 vccd1 vccd1 _6313_/D sky130_fd_sc_hd__clkbuf_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5034_ _5007_/A _5215_/B _5355_/B _5011_/A vssd1 vssd1 vccd1 vccd1 _5035_/B sky130_fd_sc_hd__a22oi_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6254__B _6254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5936_ _5936_/A _5937_/B vssd1 vssd1 vccd1 vccd1 _5936_/X sky130_fd_sc_hd__and2_1
XFILLER_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5867_ _5867_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5867_/Y sky130_fd_sc_hd__nor2_1
X_4818_ _4818_/A _4818_/B _4840_/A vssd1 vssd1 vccd1 vccd1 _4819_/B sky130_fd_sc_hd__and3_1
X_5798_ _5867_/A _5778_/A _5797_/X _3383_/A vssd1 vssd1 vccd1 vccd1 _5801_/C sky130_fd_sc_hd__a22oi_2
X_4749_ _4749_/A vssd1 vssd1 vccd1 vccd1 _4787_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3788__B _4166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4412__B _4412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3309__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3982_ _5085_/A _4168_/B _4021_/B _3981_/Y vssd1 vssd1 vccd1 vccd1 _3984_/B sky130_fd_sc_hd__a31o_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5721_ _5773_/A _5717_/Y _5815_/A _5719_/Y _5720_/Y vssd1 vssd1 vccd1 vccd1 _5744_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5652_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603_ _4603_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__xor2_1
X_5583_ _5711_/A _5630_/A vssd1 vssd1 vccd1 vccd1 _5583_/X sky130_fd_sc_hd__or2_1
X_4534_ _4534_/A _4534_/B vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__xor2_4
XANTENNA__3219__A _3220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4465_ _4328_/B _4465_/B vssd1 vssd1 vccd1 vccd1 _4465_/X sky130_fd_sc_hd__and2b_1
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4396_ _5489_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__nand2_1
X_6204_ _6352_/Q _6353_/Q _6204_/C vssd1 vssd1 vccd1 vccd1 _6204_/X sky130_fd_sc_hd__and3_1
X_3416_ _3548_/A _3416_/B vssd1 vssd1 vccd1 vccd1 _3416_/X sky130_fd_sc_hd__and2_1
XFILLER_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3347_ _3516_/A vssd1 vssd1 vccd1 vccd1 _3645_/B sky130_fd_sc_hd__clkbuf_2
X_6135_ _6325_/Q _6324_/Q _6327_/Q _6326_/Q vssd1 vssd1 vccd1 vccd1 _6135_/X sky130_fd_sc_hd__and4_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6066_ _6066_/A vssd1 vssd1 vccd1 vccd1 _6305_/D sky130_fd_sc_hd__clkbuf_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5017_ _5026_/A _5026_/B _5016_/X vssd1 vssd1 vccd1 vccd1 _5019_/B sky130_fd_sc_hd__a21oi_1
XFILLER_73_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3278_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5919_ _5919_/A vssd1 vssd1 vccd1 vccd1 _6282_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4513__A _4560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_46 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3760__A1 _3693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5265__A1 _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4250_ _4250_/A _4250_/B vssd1 vssd1 vccd1 vccd1 _4251_/B sky130_fd_sc_hd__nand2_1
X_4181_ _4181_/A _4181_/B vssd1 vssd1 vccd1 vccd1 _4472_/A sky130_fd_sc_hd__or2_2
X_3201_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3201_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3965_ _3965_/A _3965_/B vssd1 vssd1 vccd1 vccd1 _4014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3896_ _3897_/A _3897_/B vssd1 vssd1 vccd1 vccd1 _3919_/B sky130_fd_sc_hd__or2_1
XFILLER_10_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5704_ _5779_/B _5814_/C _5813_/B vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__o21ai_2
X_5635_ _5642_/A _5635_/B vssd1 vssd1 vccd1 vccd1 _5637_/B sky130_fd_sc_hd__xnor2_1
X_5566_ _5566_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _5676_/A sky130_fd_sc_hd__xnor2_2
X_4517_ _4511_/X _4515_/X _4617_/B vssd1 vssd1 vccd1 vccd1 _5746_/B sky130_fd_sc_hd__o21bai_1
X_5497_ _5497_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4448_ _5512_/A vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__clkbuf_2
X_4379_ _4403_/A _4403_/B _4378_/Y vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__a21o_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6127_/B sky130_fd_sc_hd__clkbuf_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6049_ _6036_/A _6036_/C _6042_/C _6048_/X _6036_/B vssd1 vssd1 vccd1 vccd1 _6051_/A
+ sky130_fd_sc_hd__a311oi_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5058__B _5099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3322__A _6281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3750_ _3782_/A _3782_/B vssd1 vssd1 vccd1 vccd1 _3987_/B sky130_fd_sc_hd__xnor2_2
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3681_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5130_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5420_ _5420_/A _5420_/B vssd1 vssd1 vccd1 vccd1 _5431_/A sky130_fd_sc_hd__xor2_2
XFILLER_64_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5351_ _5381_/A _5382_/B _5382_/C _5383_/A vssd1 vssd1 vccd1 vccd1 _5361_/A sky130_fd_sc_hd__and4_1
X_5282_ _5282_/A _5282_/B vssd1 vssd1 vccd1 vccd1 _5309_/A sky130_fd_sc_hd__xnor2_2
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4302_ _4303_/A _4332_/A vssd1 vssd1 vccd1 vccd1 _4317_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4233_ _4233_/A _4233_/B vssd1 vssd1 vccd1 vccd1 _4257_/A sky130_fd_sc_hd__xnor2_4
XFILLER_114_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _4164_/A _4164_/B vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _4095_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__or2_1
XFILLER_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4328__A _4465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3232__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _4997_/A _4997_/B vssd1 vssd1 vccd1 vccd1 _5559_/A sky130_fd_sc_hd__xnor2_2
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3948_ _3948_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _3949_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3879_ _5646_/A _4484_/B _3879_/C vssd1 vssd1 vccd1 vccd1 _3879_/X sky130_fd_sc_hd__and3_1
X_5618_ _5618_/A _5618_/B vssd1 vssd1 vccd1 vccd1 _5618_/Y sky130_fd_sc_hd__nand2_1
X_5549_ _5192_/X _5571_/A _5565_/B _5564_/A vssd1 vssd1 vccd1 vccd1 _5597_/B sky130_fd_sc_hd__a31o_2
XFILLER_3_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6345_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3403__B1 _4769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3317__A _3318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_616 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4920_ _4920_/A _4920_/B vssd1 vssd1 vccd1 vccd1 _4920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4851_ _4865_/A _4857_/A vssd1 vssd1 vccd1 vccd1 _4853_/B sky130_fd_sc_hd__xnor2_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ _5180_/C vssd1 vssd1 vccd1 vccd1 _3950_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__xnor2_4
X_6521_ _6521_/A _3229_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
X_3733_ _3733_/A vssd1 vssd1 vccd1 vccd1 _3734_/B sky130_fd_sc_hd__clkbuf_2
X_3664_ _3686_/A _3664_/B _3664_/C vssd1 vssd1 vccd1 vccd1 _3686_/B sky130_fd_sc_hd__nand3_1
XFILLER_9_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _5403_/A _5403_/B vssd1 vssd1 vccd1 vccd1 _5409_/B sky130_fd_sc_hd__xnor2_1
X_6383_ _6383_/CLK _6383_/D vssd1 vssd1 vccd1 vccd1 _6383_/Q sky130_fd_sc_hd__dfxtp_1
X_3595_ _3595_/A _3595_/B vssd1 vssd1 vccd1 vccd1 _3615_/A sky130_fd_sc_hd__xnor2_1
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5334_ _5334_/A _5334_/B vssd1 vssd1 vccd1 vccd1 _5360_/B sky130_fd_sc_hd__or2_1
X_5265_ _5268_/A _5263_/X _5264_/X vssd1 vssd1 vccd1 vccd1 _5578_/C sky130_fd_sc_hd__o21a_1
X_4216_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4217_/A sky130_fd_sc_hd__xnor2_1
X_5196_ _5230_/A _5196_/B _5196_/C vssd1 vssd1 vccd1 vccd1 _5198_/A sky130_fd_sc_hd__and3_1
X_4147_ _4340_/B vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_18_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4078_ _4083_/B _4078_/B vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_359 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_502 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3380_ _3380_/A _5936_/A _3380_/C vssd1 vssd1 vccd1 vccd1 _5691_/D sky130_fd_sc_hd__or3_1
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5050_/A _5050_/B vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__xor2_1
X_4001_ _4323_/A vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4606__A _4621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _6270_/A vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__buf_2
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4903_ _4898_/A _5325_/C _4764_/A _4312_/A vssd1 vssd1 vccd1 vccd1 _5289_/A sky130_fd_sc_hd__a2bb2o_1
X_5883_ _5891_/B vssd1 vssd1 vccd1 vccd1 _5899_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4834_ _4835_/A _4835_/B vssd1 vssd1 vccd1 vccd1 _4838_/B sky130_fd_sc_hd__xnor2_1
X_4765_ _4652_/A _4764_/Y _4757_/B vssd1 vssd1 vccd1 vccd1 _4783_/A sky130_fd_sc_hd__o21a_1
X_6504_ _6504_/A _3208_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_3716_ _3717_/A _3717_/C _3717_/B vssd1 vssd1 vccd1 vccd1 _3718_/C sky130_fd_sc_hd__a21o_1
XFILLER_107_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4696_ _4930_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _4698_/C sky130_fd_sc_hd__xnor2_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3647_/A _3647_/B _3647_/C vssd1 vssd1 vccd1 vccd1 _3649_/B sky130_fd_sc_hd__or3_1
XANTENNA__4343__A1 _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6366_ _6383_/CLK _6366_/D vssd1 vssd1 vccd1 vccd1 _6366_/Q sky130_fd_sc_hd__dfxtp_1
X_3578_ _3580_/C _3578_/B vssd1 vssd1 vccd1 vccd1 _3595_/B sky130_fd_sc_hd__xor2_1
XFILLER_114_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5317_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5357_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6297_ _6345_/CLK _6297_/D vssd1 vssd1 vccd1 vccd1 _6297_/Q sky130_fd_sc_hd__dfxtp_1
X_5248_ _5410_/B vssd1 vssd1 vccd1 vccd1 _5486_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5179_ _5179_/A _5179_/B _5179_/C vssd1 vssd1 vccd1 vccd1 _5186_/A sky130_fd_sc_hd__nand3_2
XFILLER_68_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4516__A _4516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4235__B _4235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5822__A1_N _5698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4550_/A _4550_/B vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__or2_1
X_4481_ _4521_/A _4495_/A _4494_/B vssd1 vssd1 vccd1 vccd1 _4492_/B sky130_fd_sc_hd__or3_1
X_3501_ _6040_/A _3653_/B _4768_/C vssd1 vssd1 vccd1 vccd1 _3697_/C sky130_fd_sc_hd__nor3_2
XFILLER_7_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3432_ _3432_/A _3432_/B vssd1 vssd1 vccd1 vccd1 _3473_/B sky130_fd_sc_hd__xnor2_1
X_6220_ _6270_/A vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__clkbuf_2
X_3363_ _4864_/B vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__clkbuf_2
X_6151_ _6337_/Q _6165_/B vssd1 vssd1 vccd1 vccd1 _6152_/A sky130_fd_sc_hd__and2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5102_ _5108_/A _5101_/B _3950_/A _5059_/B vssd1 vssd1 vccd1 vccd1 _5104_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6359_/Q _6096_/B vssd1 vssd1 vccd1 vccd1 _6083_/A sky130_fd_sc_hd__and2_1
X_3294_ _3294_/A vssd1 vssd1 vccd1 vccd1 _3294_/Y sky130_fd_sc_hd__inv_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5196_/B vssd1 vssd1 vccd1 vccd1 _5355_/B sky130_fd_sc_hd__buf_2
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5935_ _5935_/A _5941_/A vssd1 vssd1 vccd1 vccd1 _5937_/B sky130_fd_sc_hd__xor2_1
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5866_ _5866_/A _5867_/B vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__and2_1
X_4817_ _4818_/B _4840_/A _4818_/A vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5167__A _5382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5797_ _5769_/X _5749_/Y _5771_/Y _5747_/X vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__a22o_1
X_4748_ _4787_/B vssd1 vssd1 vccd1 vccd1 _4879_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4679_ _4722_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4682_/C sky130_fd_sc_hd__or2b_1
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6349_ _6357_/CLK _6349_/D vssd1 vssd1 vccd1 vccd1 _6349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5630__A _5630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4246__A _6280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5761__A1_N _5901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3981_ _3981_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _3981_/Y sky130_fd_sc_hd__nor2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _5714_/A _5699_/B _5777_/A vssd1 vssd1 vccd1 vccd1 _5720_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6529__48 vssd1 vssd1 vccd1 vccd1 _6529__48/HI _6529_/A sky130_fd_sc_hd__conb_1
XANTENNA__4603__B _4603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5651_ _5865_/A _5651_/B _5651_/C vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__or3_1
X_5582_ _5582_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5630_/A sky130_fd_sc_hd__xnor2_4
X_4602_ _4621_/B _4606_/B vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4533_ _4603_/A vssd1 vssd1 vccd1 vccd1 _5735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4464_ _4534_/A _4534_/B _4463_/Y vssd1 vssd1 vccd1 vccd1 _4538_/B sky130_fd_sc_hd__a21o_1
X_6203_ _6356_/Q _6355_/Q _6358_/Q _6357_/Q vssd1 vssd1 vccd1 vccd1 _6204_/C sky130_fd_sc_hd__and4_1
XANTENNA__3235__A _3239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4395_ _4397_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__xnor2_1
X_3415_ _3548_/A _3416_/B vssd1 vssd1 vccd1 vccd1 _3469_/B sky130_fd_sc_hd__xor2_1
XFILLER_112_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6134_ _6329_/Q _6328_/Q _6331_/Q _6330_/Q vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__and4_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _6287_/Q vssd1 vssd1 vccd1 vccd1 _3516_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _6140_/A input5/X vssd1 vssd1 vccd1 vccd1 _6066_/A sky130_fd_sc_hd__and2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__buf_8
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5016_ _5015_/B _5016_/B vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__and2b_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5544__A_N _5308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5918_ _6332_/Q _5980_/B vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__and2_1
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4513__B _4626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5849_ _5844_/X _5847_/X _5848_/X vssd1 vssd1 vccd1 vccd1 _5849_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4796__D _4796_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4180_ _4180_/A _4180_/B _4180_/C vssd1 vssd1 vccd1 vccd1 _4181_/B sky130_fd_sc_hd__nor3_1
X_3200_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3200_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3964_ _3964_/A _3964_/B vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__or2_1
XANTENNA__5964__B1 _5952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3895_ _3895_/A _3900_/A vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__xor2_1
XFILLER_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5703_ _5703_/A _5759_/A vssd1 vssd1 vccd1 vccd1 _5703_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5716__B1 _5724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5634_ _5634_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5639_/A sky130_fd_sc_hd__xnor2_1
X_5565_ _5571_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _5566_/B sky130_fd_sc_hd__nand2_1
X_4516_ _4516_/A _4516_/B vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__xnor2_1
X_5496_ _5426_/A _5489_/B _5490_/A _5488_/A vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__a31o_1
XFILLER_2_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4447_ _5485_/A vssd1 vssd1 vccd1 vccd1 _5512_/A sky130_fd_sc_hd__inv_2
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input6_A io_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ _4378_/A _4378_/B vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__nor2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6189_/B vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3329_ _4929_/A vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6048_ _6040_/A _6300_/Q _6046_/B vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__o21a_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5355__A _5355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5249__B _5486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3680_ _5294_/A vssd1 vssd1 vccd1 vccd1 _5165_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5350_ _5410_/A _5469_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5383_/A sky130_fd_sc_hd__and3_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5281_ _5281_/A _5281_/B vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4301_ _5411_/A _4301_/B vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _4059_/A _4235_/B _4234_/B _4231_/X vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__a31o_2
X_4163_ _4182_/A _4182_/B vssd1 vssd1 vccd1 vccd1 _4164_/B sky130_fd_sc_hd__and2b_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4106_/B sky130_fd_sc_hd__inv_2
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _4996_/A _4996_/B vssd1 vssd1 vccd1 vccd1 _4997_/B sky130_fd_sc_hd__xnor2_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3947_ _5064_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4063__B _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3878_ _3906_/B vssd1 vssd1 vccd1 vccd1 _4484_/B sky130_fd_sc_hd__clkbuf_2
X_6597_ _6597_/A _3315_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_5617_ _5698_/A _5619_/B _5616_/Y vssd1 vssd1 vccd1 vccd1 _5618_/B sky130_fd_sc_hd__a21o_1
X_5548_ _5189_/Y _5546_/A _5154_/B _5156_/X vssd1 vssd1 vccd1 vccd1 _5564_/A sky130_fd_sc_hd__o211a_1
XFILLER_3_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6513__32 vssd1 vssd1 vccd1 vccd1 _6513__32/HI _6513_/A sky130_fd_sc_hd__conb_1
X_5479_ _5482_/A _5482_/B vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__or2b_1
XANTENNA__4519__A _5710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4979__A1 _5627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5085__A _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4754__A1_N _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3987__B _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4850_ _4856_/A _4850_/B vssd1 vssd1 vccd1 vccd1 _4857_/A sky130_fd_sc_hd__xor2_1
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ _4079_/A vssd1 vssd1 vccd1 vccd1 _5180_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _4920_/A _4920_/B vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__xor2_4
X_6520_ _6520_/A _3228_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_3732_ _3377_/A _3733_/A _3734_/C vssd1 vssd1 vccd1 vccd1 _3735_/A sky130_fd_sc_hd__a21o_1
XFILLER_9_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3663_ _3663_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3664_/C sky130_fd_sc_hd__or2_1
X_5402_ _5420_/A _5420_/B _5401_/X vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__o21a_1
X_6382_ _6383_/CLK _6382_/D vssd1 vssd1 vccd1 vccd1 _6382_/Q sky130_fd_sc_hd__dfxtp_1
X_5333_ _5332_/B _5333_/B vssd1 vssd1 vccd1 vccd1 _5334_/B sky130_fd_sc_hd__and2b_1
X_3594_ _3594_/A _3594_/B vssd1 vssd1 vccd1 vccd1 _3595_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5264_ _5264_/A _5264_/B _5267_/B vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__or3_1
X_4215_ _4233_/A _4233_/B _4214_/X vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__a21oi_2
X_5195_ _5195_/A _5273_/B vssd1 vssd1 vccd1 vccd1 _5196_/C sky130_fd_sc_hd__and2_1
XANTENNA__5442__B _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ _5246_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3243__A _3245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4077_ _4075_/A _4075_/B _4108_/A vssd1 vssd1 vccd1 vccd1 _4078_/B sky130_fd_sc_hd__o21ba_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4979_ _5627_/A _4994_/B _4978_/C vssd1 vssd1 vccd1 vccd1 _4980_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3328__A _5011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ _5276_/A vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5951_ _5951_/A _5951_/B _5951_/C vssd1 vssd1 vccd1 vccd1 _5951_/X sky130_fd_sc_hd__and3_1
X_4902_ _4902_/A _4902_/B vssd1 vssd1 vccd1 vccd1 _5247_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5882_ _5879_/A _5879_/B _5876_/A vssd1 vssd1 vccd1 vccd1 _5886_/A sky130_fd_sc_hd__o21ai_1
X_4833_ _4833_/A _4855_/A vssd1 vssd1 vccd1 vccd1 _4835_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5368__A1 _5246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4764_ _4764_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4764_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6503_ _6503_/A _3207_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_3715_ _3715_/A _3715_/B vssd1 vssd1 vccd1 vccd1 _3717_/B sky130_fd_sc_hd__nor2_1
X_4695_ _4950_/B _4695_/B vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3238__A _3239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _3696_/A _3600_/B _3645_/D _3645_/B vssd1 vssd1 vccd1 vccd1 _3647_/C sky130_fd_sc_hd__a22oi_2
X_6365_ _6375_/CLK _6365_/D vssd1 vssd1 vccd1 vccd1 _6365_/Q sky130_fd_sc_hd__dfxtp_1
X_3577_ _3580_/A _4882_/A vssd1 vssd1 vccd1 vccd1 _3578_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5316_ _5358_/A _5316_/B vssd1 vssd1 vccd1 vccd1 _5341_/B sky130_fd_sc_hd__nand2_1
X_6296_ _6335_/CLK _6296_/D vssd1 vssd1 vccd1 vccd1 _6296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5172__B _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5247_ _5247_/A _5290_/A vssd1 vssd1 vccd1 vccd1 _5410_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5178_ _5176_/A _5176_/B _5214_/A vssd1 vssd1 vccd1 vccd1 _5179_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4129_ _5098_/A _4168_/B _4120_/X _4124_/B vssd1 vssd1 vccd1 vccd1 _4137_/A sky130_fd_sc_hd__a31o_1
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3420__B _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3790__B1 _3947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6589__105 vssd1 vssd1 vccd1 vccd1 _6589__105/HI _6589_/A sky130_fd_sc_hd__conb_1
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3500_ _3642_/B _3499_/C _3476_/Y vssd1 vssd1 vccd1 vccd1 _3508_/B sky130_fd_sc_hd__a21boi_1
XFILLER_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _4537_/A _4536_/A _4536_/B _4521_/B _4017_/A vssd1 vssd1 vccd1 vccd1 _4494_/B
+ sky130_fd_sc_hd__a311oi_2
XFILLER_7_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3431_ _4842_/B _3692_/B vssd1 vssd1 vccd1 vccd1 _3432_/B sky130_fd_sc_hd__nand2_1
X_6150_ _6150_/A vssd1 vssd1 vccd1 vccd1 _6337_/D sky130_fd_sc_hd__clkbuf_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _6284_/Q vssd1 vssd1 vccd1 vccd1 _4864_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5101_ _5108_/A _5101_/B _5180_/C _5059_/B vssd1 vssd1 vccd1 vccd1 _5104_/A sky130_fd_sc_hd__or4bb_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3294_/A vssd1 vssd1 vccd1 vccd1 _3293_/Y sky130_fd_sc_hd__inv_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A vssd1 vssd1 vccd1 vccd1 _6312_/D sky130_fd_sc_hd__clkbuf_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/A _5070_/A vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__nor2_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5934_ _5924_/X _5926_/X _5927_/X _5925_/Y vssd1 vssd1 vccd1 vccd1 _5941_/A sky130_fd_sc_hd__o22a_1
X_5865_ _5865_/A _5877_/A vssd1 vssd1 vccd1 vccd1 _5867_/B sky130_fd_sc_hd__xnor2_1
X_4816_ _4818_/B _4816_/B _4816_/C vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5796_ _6368_/Q vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4747_ _4747_/A _4747_/B vssd1 vssd1 vccd1 vccd1 _4920_/A sky130_fd_sc_hd__xor2_4
X_6555__71 vssd1 vssd1 vccd1 vccd1 _6555__71/HI _6555_/A sky130_fd_sc_hd__conb_1
XFILLER_107_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4678_ _4645_/Y _4712_/A _4682_/B vssd1 vssd1 vccd1 vccd1 _4722_/B sky130_fd_sc_hd__a21boi_1
XFILLER_107_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5513__B2 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3629_ _3629_/A _3629_/B vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6348_ _6357_/CLK _6348_/D vssd1 vssd1 vccd1 vccd1 _6348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6279_ _6359_/CLK _6279_/D vssd1 vssd1 vccd1 vccd1 _6279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4527__A _4560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_46 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_528 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ _3981_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__xor2_1
XFILLER_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5268__A _5268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5650_ _5511_/B _5610_/B _4138_/A vssd1 vssd1 vccd1 vccd1 _5651_/C sky130_fd_sc_hd__a21bo_1
XFILLER_15_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4601_ _4550_/X _4556_/Y _4562_/Y _4563_/Y _4600_/X vssd1 vssd1 vccd1 vccd1 _4611_/A
+ sky130_fd_sc_hd__o221a_1
X_5581_ _5703_/A _5672_/A vssd1 vssd1 vccd1 vccd1 _5581_/X sky130_fd_sc_hd__xor2_1
X_4532_ _4532_/A _4532_/B vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__xnor2_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4463_ _4463_/A _4463_/B vssd1 vssd1 vccd1 vccd1 _4463_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5715__B _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3506__B1 _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6202_ _6202_/A vssd1 vssd1 vccd1 vccd1 _6358_/D sky130_fd_sc_hd__clkbuf_1
X_3414_ _6289_/Q _3436_/A _3436_/B vssd1 vssd1 vccd1 vccd1 _3416_/B sky130_fd_sc_hd__and3_1
X_4394_ _5416_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4397_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6133_ _6133_/A vssd1 vssd1 vccd1 vccd1 _6331_/D sky130_fd_sc_hd__clkbuf_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _5935_/A vssd1 vssd1 vccd1 vccd1 _3381_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3276_ _3276_/A vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6064_ _6254_/B _6064_/B vssd1 vssd1 vccd1 vccd1 _6304_/D sky130_fd_sc_hd__nor2_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5016_/B _5015_/B vssd1 vssd1 vccd1 vccd1 _5026_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5450__B _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3251__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5917_ _5917_/A vssd1 vssd1 vccd1 vccd1 _6281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _6381_/Q _5846_/X _5822_/X _6382_/Q vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5734__B2 _5733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5779_ _5779_/A _5779_/B _6302_/Q vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__or3_2
XANTENNA__5906__A _5906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3963_ _4010_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _3964_/B sky130_fd_sc_hd__and2b_1
X_3894_ _3901_/A _3894_/B vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__xor2_1
X_5702_ _5702_/A _5757_/A vssd1 vssd1 vccd1 vccd1 _5702_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5633_ _5633_/A _5633_/B vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__or2_1
X_5564_ _5564_/A _5192_/X vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__or2b_1
XFILLER_12_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4515_ _4618_/A _4618_/B vssd1 vssd1 vccd1 vccd1 _4515_/X sky130_fd_sc_hd__and2_1
X_5495_ _5497_/A _5497_/B vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__and2b_1
X_4446_ _5514_/A _4449_/B _4445_/Y vssd1 vssd1 vccd1 vccd1 _4451_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4152__B1 _4153_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4377_ _4377_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4403_/B sky130_fd_sc_hd__xnor2_1
X_3328_ _5011_/A vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A vssd1 vssd1 vccd1 vccd1 _6324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3259_ _3263_/A vssd1 vssd1 vccd1 vccd1 _3259_/Y sky130_fd_sc_hd__inv_2
X_6047_ _6055_/A _6047_/B vssd1 vssd1 vccd1 vccd1 _6050_/A sky130_fd_sc_hd__and2_1
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__B _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4540__A _5724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5636__A _5637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5355__B _5355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4153__C _4153_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5280_ _5277_/A _5277_/B _5279_/Y vssd1 vssd1 vccd1 vccd1 _5310_/A sky130_fd_sc_hd__o21ba_2
X_4300_ _6278_/Q vssd1 vssd1 vccd1 vccd1 _5411_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _4226_/Y _4229_/X _5314_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4162_ _4162_/A _4162_/B vssd1 vssd1 vccd1 vccd1 _4182_/B sky130_fd_sc_hd__xnor2_2
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4093_ _4093_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4995_ _4993_/Y _4989_/A _4995_/S vssd1 vssd1 vccd1 vccd1 _4996_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3946_ _3944_/A _3944_/B _3945_/X vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__o21ba_1
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3877_ _3877_/A vssd1 vssd1 vccd1 vccd1 _5646_/A sky130_fd_sc_hd__buf_2
XFILLER_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6596_ _6596_/A _3316_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_5616_ _5672_/A _5616_/B vssd1 vssd1 vccd1 vccd1 _5616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547_ _5579_/A _5570_/B _5571_/B vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__a21bo_1
X_5478_ _5478_/A _5478_/B vssd1 vssd1 vccd1 vccd1 _5482_/B sky130_fd_sc_hd__xor2_1
X_4429_ _5471_/A _4430_/B vssd1 vssd1 vccd1 vccd1 _4429_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3800_ _5199_/A vssd1 vssd1 vccd1 vccd1 _4079_/A sky130_fd_sc_hd__clkbuf_2
X_4780_ _4782_/A _4782_/B _4779_/X vssd1 vssd1 vccd1 vccd1 _4920_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3731_ _3731_/A _3731_/B vssd1 vssd1 vccd1 vccd1 _3759_/B sky130_fd_sc_hd__nand2_1
X_3662_ _4644_/A _3644_/B _3495_/B _3505_/A _3502_/X vssd1 vssd1 vccd1 vccd1 _3663_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5401_ _5401_/A _5401_/B vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__or2_1
X_6381_ _6383_/CLK _6381_/D vssd1 vssd1 vccd1 vccd1 _6381_/Q sky130_fd_sc_hd__dfxtp_1
X_3593_ _3599_/A _3598_/B _3592_/X vssd1 vssd1 vccd1 vccd1 _3615_/B sky130_fd_sc_hd__a21oi_1
X_5332_ _5333_/B _5332_/B vssd1 vssd1 vccd1 vccd1 _5334_/A sky130_fd_sc_hd__and2b_1
XFILLER_102_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5263_ _5267_/A _5267_/B vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__and2b_1
X_4214_ _4206_/B _4214_/B vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__and2b_1
X_5194_ _5177_/A _5177_/B _5177_/C vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5442__C _5471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _4145_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__and2_1
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4076_ _4115_/A _4076_/B _4076_/C vssd1 vssd1 vccd1 vccd1 _4108_/A sky130_fd_sc_hd__and3_1
XFILLER_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4074__B _4396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4978_ _4978_/A _4994_/B _4978_/C vssd1 vssd1 vccd1 vccd1 _4988_/B sky130_fd_sc_hd__and3_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3929_ _4486_/A _3929_/B vssd1 vssd1 vccd1 vccd1 _3931_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6579_ _6579_/A _3293_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
XFILLER_3_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4249__B _4250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5950_ _5940_/A _3381_/B _5937_/A _5949_/X vssd1 vssd1 vccd1 vccd1 _5951_/C sky130_fd_sc_hd__o31ai_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4901_ _4908_/A _4908_/B _4908_/C vssd1 vssd1 vccd1 vccd1 _5203_/B sky130_fd_sc_hd__a21o_1
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5881_ _5733_/X _5857_/X _5880_/Y _5872_/X vssd1 vssd1 vccd1 vccd1 _6276_/D sky130_fd_sc_hd__o211a_1
X_4832_ _4833_/A _4832_/B _4832_/C vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__nand3_1
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__xnor2_1
X_6502_ _6502_/A _3206_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_3714_ _3713_/B _3714_/B vssd1 vssd1 vccd1 vccd1 _3715_/B sky130_fd_sc_hd__and2b_1
X_4694_ _4694_/A _4694_/B _4694_/C vssd1 vssd1 vccd1 vccd1 _4695_/B sky130_fd_sc_hd__and3_1
X_3645_ _3696_/A _3645_/B _3645_/C _3645_/D vssd1 vssd1 vccd1 vccd1 _3647_/B sky130_fd_sc_hd__and4_1
XFILLER_20_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6364_ _6375_/CLK _6364_/D vssd1 vssd1 vccd1 vccd1 _6364_/Q sky130_fd_sc_hd__dfxtp_1
X_3576_ _3576_/A vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__clkbuf_2
X_5315_ _5315_/A _5315_/B vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__xor2_2
X_6295_ _6335_/CLK _6295_/D vssd1 vssd1 vccd1 vccd1 _6295_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3254__A _3257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5246_ _5246_/A _5246_/B vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _5177_/A _5177_/B _5177_/C vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__and3_1
XFILLER_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _5236_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4059_ _4059_/A vssd1 vssd1 vccd1 vccd1 _5183_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3790__A1 _5011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4707__B _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5819__A _5819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3339__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3430_ _3592_/A vssd1 vssd1 vccd1 vccd1 _4842_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_112_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5273__B _5273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3361_ _4692_/A vssd1 vssd1 vccd1 vccd1 _3380_/A sky130_fd_sc_hd__buf_2
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5100_ _5098_/A _5236_/B _5098_/C vssd1 vssd1 vccd1 vccd1 _5101_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3505__C _3505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6080_ _6311_/Q _6096_/B vssd1 vssd1 vccd1 vccd1 _6081_/A sky130_fd_sc_hd__and2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5031_ _5091_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__nand2_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3294_/A vssd1 vssd1 vccd1 vccd1 _3292_/Y sky130_fd_sc_hd__inv_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _5937_/A _5930_/X _5932_/Y vssd1 vssd1 vccd1 vccd1 _6284_/D sky130_fd_sc_hd__a21oi_1
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5864_ _5851_/X _5853_/X _5854_/X _5852_/Y vssd1 vssd1 vccd1 vccd1 _5877_/A sky130_fd_sc_hd__o22a_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4549__B1 _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4815_ _4815_/A _4877_/C vssd1 vssd1 vccd1 vccd1 _4816_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3249__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5795_ _5741_/A _5778_/X _5794_/X _5694_/X vssd1 vssd1 vccd1 vccd1 _5795_/X sky130_fd_sc_hd__o2bb2a_1
X_4746_ _4746_/A _4746_/B vssd1 vssd1 vccd1 vccd1 _4926_/A sky130_fd_sc_hd__nor2_2
XFILLER_31_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4677_ _4677_/A _4677_/B vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__xnor2_1
X_3628_ _3627_/A _3627_/B _3627_/C vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__a21o_1
X_6347_ _6357_/CLK _6347_/D vssd1 vssd1 vccd1 vccd1 _6347_/Q sky130_fd_sc_hd__dfxtp_1
X_6570__86 vssd1 vssd1 vccd1 vccd1 _6570__86/HI _6570_/A sky130_fd_sc_hd__conb_1
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3559_ _4787_/A _3559_/B _3580_/C vssd1 vssd1 vccd1 vccd1 _3560_/C sky130_fd_sc_hd__and3_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6278_ _6359_/CLK _6278_/D vssd1 vssd1 vccd1 vccd1 _6278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5229_ _5224_/A _5225_/X _5216_/X _5221_/B vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__a211oi_1
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4527__B _4626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5358__B _5358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4262__B _4340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4600_ _4562_/Y _4563_/Y _4564_/Y _4571_/Y _4599_/X vssd1 vssd1 vccd1 vccd1 _4600_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5580_ _5580_/A _5580_/B vssd1 vssd1 vccd1 vccd1 _5672_/A sky130_fd_sc_hd__xnor2_4
X_4531_ _4531_/A _4531_/B vssd1 vssd1 vccd1 vccd1 _4532_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4462_ _4593_/A _4593_/B _4461_/X vssd1 vssd1 vccd1 vccd1 _4534_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6201_ _6357_/Q _6201_/B vssd1 vssd1 vccd1 vccd1 _6202_/A sky130_fd_sc_hd__and2_1
X_3413_ _3386_/A _3406_/X _6295_/Q _3517_/A vssd1 vssd1 vccd1 vccd1 _3436_/B sky130_fd_sc_hd__a22oi_2
X_4393_ _4393_/A _4417_/A vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__nor2_1
X_3344_ _4898_/A vssd1 vssd1 vccd1 vccd1 _5935_/A sky130_fd_sc_hd__clkbuf_2
X_6132_ _6330_/Q _6146_/B vssd1 vssd1 vccd1 vccd1 _6133_/A sky130_fd_sc_hd__and2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4628__A _4796_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3275_ _3276_/A vssd1 vssd1 vccd1 vccd1 _3275_/Y sky130_fd_sc_hd__inv_2
X_6063_ _6063_/A _6063_/B vssd1 vssd1 vccd1 vccd1 _6064_/B sky130_fd_sc_hd__xor2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5012_/A _5032_/A _5028_/A vssd1 vssd1 vccd1 vccd1 _5015_/B sky130_fd_sc_hd__o21ba_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_587 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5916_ _5914_/X _5916_/B vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__and2b_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5847_ _6380_/Q _5825_/Y _5846_/X _6381_/Q vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5778_ _5778_/A vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4729_ _4879_/C vssd1 vssd1 vccd1 vccd1 _4877_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4170__A1 _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6534__53 vssd1 vssd1 vccd1 vccd1 _6534__53/HI _6534_/A sky130_fd_sc_hd__conb_1
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3962_ _3877_/A _4063_/B _3956_/B _3961_/Y vssd1 vssd1 vccd1 vccd1 _4010_/B sky130_fd_sc_hd__a31o_1
XFILLER_90_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5701_ _5779_/A _5701_/B _5814_/C vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__or3_2
XFILLER_50_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3893_ _3916_/A _3893_/B vssd1 vssd1 vccd1 vccd1 _3894_/B sky130_fd_sc_hd__and2_1
XFILLER_50_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5632_ _5629_/A _5630_/A _5629_/B _5631_/Y vssd1 vssd1 vccd1 vccd1 _5633_/B sky130_fd_sc_hd__o31a_1
X_5563_ _5711_/A vssd1 vssd1 vccd1 vccd1 _5683_/B sky130_fd_sc_hd__inv_2
X_4514_ _4555_/A _5702_/A vssd1 vssd1 vccd1 vccd1 _4618_/B sky130_fd_sc_hd__xnor2_1
X_5494_ _5501_/A _5501_/B vssd1 vssd1 vccd1 vccd1 _5497_/B sky130_fd_sc_hd__and2_1
X_4445_ _4445_/A _4587_/A vssd1 vssd1 vccd1 vccd1 _4445_/Y sky130_fd_sc_hd__nor2_1
X_6540__56 vssd1 vssd1 vccd1 vccd1 _6540__56/HI _6540_/A sky130_fd_sc_hd__conb_1
X_4376_ _5489_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3327_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__clkbuf_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6140_/A input3/X vssd1 vssd1 vccd1 vccd1 _6116_/A sky130_fd_sc_hd__and2_1
XANTENNA__3262__A _3263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3258_ _3258_/A vssd1 vssd1 vccd1 vccd1 _3263_/A sky130_fd_sc_hd__buf_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6061_/B _6046_/B vssd1 vssd1 vccd1 vccd1 _6047_/B sky130_fd_sc_hd__or2_1
X_3189_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4540__B _4583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5099__A _5099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4450__B _5511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4230_ _5314_/A _3940_/B _4226_/Y _4229_/X vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__a211o_1
X_4161_ _4168_/C _4161_/B vssd1 vssd1 vccd1 vccd1 _4182_/A sky130_fd_sc_hd__xor2_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4092_ _4098_/C _4092_/B vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4994_ _5605_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _4995_/S sky130_fd_sc_hd__nand2_1
X_3945_ _5064_/A _4235_/B _3972_/B vssd1 vssd1 vccd1 vccd1 _3945_/X sky130_fd_sc_hd__and3_1
XFILLER_23_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5737__A _5737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3876_ _3881_/A _3881_/B vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__nand2_1
X_5615_ _5672_/A _5616_/B vssd1 vssd1 vccd1 vccd1 _5619_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3257__A _3257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6595_ _6595_/A _3319_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_5546_ _5546_/A _5546_/B _5546_/C vssd1 vssd1 vccd1 vccd1 _5571_/B sky130_fd_sc_hd__or3_1
X_5477_ _5472_/A _5472_/B _5476_/X vssd1 vssd1 vccd1 vccd1 _5482_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4428_ _6274_/Q vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4359_ _5411_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _6031_/B vssd1 vssd1 vccd1 vccd1 _6046_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5625__A1 _5755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6504__23 vssd1 vssd1 vccd1 vccd1 _6504__23/HI _6504_/A sky130_fd_sc_hd__conb_1
XFILLER_89_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5813__C _6060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4726__A _4726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3730_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3758_/A sky130_fd_sc_hd__or2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ _3661_/A _3807_/B _3661_/C vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__and3_1
X_5400_ _5401_/A _5401_/B vssd1 vssd1 vccd1 vccd1 _5420_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3592_ _3592_/A _6284_/Q _3645_/C _3696_/B vssd1 vssd1 vccd1 vccd1 _3592_/X sky130_fd_sc_hd__and4_1
X_6380_ _6383_/CLK _6380_/D vssd1 vssd1 vccd1 vccd1 _6380_/Q sky130_fd_sc_hd__dfxtp_1
X_5331_ _5329_/A _5329_/B _5370_/A vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__o21bai_1
XFILLER_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5262_ _5237_/Y _5241_/X _5282_/B _5261_/Y vssd1 vssd1 vccd1 vccd1 _5267_/B sky130_fd_sc_hd__o31a_1
X_4213_ _4213_/A _4213_/B vssd1 vssd1 vccd1 vccd1 _4233_/B sky130_fd_sc_hd__xor2_4
XFILLER_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5193_ _5189_/Y _5190_/X _5183_/C _5186_/B vssd1 vssd1 vccd1 vccd1 _5546_/B sky130_fd_sc_hd__o211a_1
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4144_ _4124_/B _4124_/C _4124_/A vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__o21ai_1
XFILLER_18_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4075_ _4075_/A _4075_/B vssd1 vssd1 vccd1 vccd1 _4076_/C sky130_fd_sc_hd__xor2_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4977_ _4988_/A _4977_/B vssd1 vssd1 vccd1 vccd1 _4978_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4594__A1 _4370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ _3928_/A _3928_/B _3928_/C vssd1 vssd1 vccd1 vccd1 _3929_/B sky130_fd_sc_hd__nor3_1
X_3859_ _4960_/A _4166_/B _3790_/X _3885_/C _3754_/B vssd1 vssd1 vccd1 vccd1 _3883_/A
+ sky130_fd_sc_hd__a32oi_2
X_6578_ _6578_/A _3291_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
XFILLER_105_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5529_ _5529_/A _5500_/A vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__or2b_1
XFILLER_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4546__A _4546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6576__92 vssd1 vssd1 vccd1 vccd1 _6576__92/HI _6576_/A sky130_fd_sc_hd__conb_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4902_/A _4902_/B vssd1 vssd1 vccd1 vccd1 _4908_/C sky130_fd_sc_hd__nand2_1
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5880_ _5910_/A _5880_/B vssd1 vssd1 vccd1 vccd1 _5880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4831_ _4829_/A _4829_/B _4852_/C vssd1 vssd1 vccd1 vccd1 _4832_/C sky130_fd_sc_hd__a21o_1
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5287__A _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4762_ _4762_/A _4797_/A vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__xnor2_2
X_3713_ _3714_/B _3713_/B vssd1 vssd1 vccd1 vccd1 _3715_/A sky130_fd_sc_hd__and2b_1
X_4693_ _4693_/A vssd1 vssd1 vccd1 vccd1 _4694_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6501_ _6501_/A _3205_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_3644_ _4651_/A _3644_/B vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6363_ _6383_/CLK _6363_/D vssd1 vssd1 vccd1 vccd1 _6363_/Q sky130_fd_sc_hd__dfxtp_1
X_3575_ _3601_/A _3644_/B _3575_/C vssd1 vssd1 vccd1 vccd1 _3594_/B sky130_fd_sc_hd__nand3_1
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5314_ _5314_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5315_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6495__14 vssd1 vssd1 vccd1 vccd1 _6495__14/HI _6495_/A sky130_fd_sc_hd__conb_1
X_6294_ _6335_/CLK _6294_/D vssd1 vssd1 vccd1 vccd1 _6294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5245_ _5245_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5257_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5176_ _5176_/A _5176_/B vssd1 vssd1 vccd1 vccd1 _5177_/C sky130_fd_sc_hd__xor2_1
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4127_ _4134_/B _4127_/B vssd1 vssd1 vccd1 vccd1 _4143_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3270__A _3270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4058_ _4041_/X _4056_/Y _4057_/X _4009_/B vssd1 vssd1 vccd1 vccd1 _4066_/A sky130_fd_sc_hd__o211a_1
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3790__A2 _4235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6295__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3355__A _4726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _4731_/A vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3294_/A vssd1 vssd1 vccd1 vccd1 _3291_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5030_ _5196_/B vssd1 vssd1 vccd1 vccd1 _5358_/B sky130_fd_sc_hd__clkbuf_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_608 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _5937_/A _5970_/A _5861_/X vssd1 vssd1 vccd1 vccd1 _5932_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5863_ _5867_/A _5857_/X _5862_/Y vssd1 vssd1 vccd1 vccd1 _6274_/D sky130_fd_sc_hd__a21oi_1
X_4814_ _4814_/A _4814_/B _4814_/C _4707_/A vssd1 vssd1 vccd1 vccd1 _4816_/B sky130_fd_sc_hd__or4b_1
XFILLER_33_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5794_ _5690_/A _5792_/X _5815_/B _5793_/X vssd1 vssd1 vccd1 vccd1 _5794_/X sky130_fd_sc_hd__o22a_1
X_4745_ _4745_/A _4745_/B _4745_/C vssd1 vssd1 vccd1 vccd1 _4746_/B sky130_fd_sc_hd__nor3_1
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5745__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4676_ _4645_/Y _4674_/X _4712_/A vssd1 vssd1 vccd1 vccd1 _4682_/B sky130_fd_sc_hd__a21o_1
X_3627_ _3627_/A _3627_/B _3627_/C vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__nand3_1
X_6346_ _6357_/CLK _6346_/D vssd1 vssd1 vccd1 vccd1 _6346_/Q sky130_fd_sc_hd__dfxtp_1
X_3558_ _4865_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _3580_/C sky130_fd_sc_hd__xnor2_2
XFILLER_103_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6277_ _6359_/CLK _6277_/D vssd1 vssd1 vccd1 vccd1 _6277_/Q sky130_fd_sc_hd__dfxtp_1
X_3489_ _3489_/A _3643_/B _3489_/C vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__nand3_1
X_5228_ _5546_/A _5546_/B _5546_/C vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__o21ai_1
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5159_ _5159_/A _5159_/B vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6595__111 vssd1 vssd1 vccd1 vccd1 _6595__111/HI _6595_/A sky130_fd_sc_hd__conb_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6546__62 vssd1 vssd1 vccd1 vccd1 _6546__62/HI _6546_/A sky130_fd_sc_hd__conb_1
XFILLER_4_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4530_ _4506_/A _4506_/B _4477_/X vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__a21o_1
XANTENNA__4951__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4461_ _4383_/B _4461_/B vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6200_ _6200_/A vssd1 vssd1 vccd1 vccd1 _6357_/D sky130_fd_sc_hd__clkbuf_1
X_3412_ _3405_/X _3406_/X _6295_/Q _3517_/A vssd1 vssd1 vccd1 vccd1 _3436_/A sky130_fd_sc_hd__a211o_1
XFILLER_98_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4392_ _5382_/A _4430_/B _4392_/C vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__and3_1
X_6131_ _6131_/A vssd1 vssd1 vccd1 vccd1 _6330_/D sky130_fd_sc_hd__clkbuf_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3343_ _3505_/A vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3276_/A vssd1 vssd1 vccd1 vccd1 _3274_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6062_ _6060_/X _6061_/X _5989_/A vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__a21bo_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5013_/A _5013_/B _5013_/C vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__and3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6208__B2 _5861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5915_ _5868_/A _5912_/X _5913_/Y _3333_/X vssd1 vssd1 vccd1 vccd1 _5916_/B sky130_fd_sc_hd__a31o_1
X_5846_ _5755_/A _5820_/X _5845_/X _5694_/X vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__o2bb2a_1
X_5777_ _5777_/A _5777_/B vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__or2_1
X_4728_ _3387_/A _5685_/A _5993_/A vssd1 vssd1 vccd1 vccd1 _4879_/C sky130_fd_sc_hd__a21o_1
X_4659_ _4659_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__xnor2_1
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6329_ _6345_/CLK _6329_/D vssd1 vssd1 vccd1 vccd1 _6329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4554__A _4555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4183__B _4337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ _3993_/A _3961_/B vssd1 vssd1 vccd1 vccd1 _3961_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5700_ _5741_/B vssd1 vssd1 vccd1 vccd1 _5700_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3892_ _3892_/A _3892_/B _3892_/C vssd1 vssd1 vccd1 vccd1 _3893_/B sky130_fd_sc_hd__or3_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5631_ _5899_/A _5634_/B vssd1 vssd1 vccd1 vccd1 _5631_/Y sky130_fd_sc_hd__nand2_1
X_5562_ _5562_/A _5562_/B vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__xnor2_4
X_4513_ _4560_/A _4626_/A vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5493_ _5493_/A _5493_/B vssd1 vssd1 vccd1 vccd1 _5501_/B sky130_fd_sc_hd__nor2_1
X_4444_ _4445_/A _4587_/A _4443_/X vssd1 vssd1 vccd1 vccd1 _4449_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4152__A2 _4412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4375_ _4378_/A _4378_/B vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__xor2_1
X_3326_ _5166_/A vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _6318_/Q _6316_/D _6110_/X _6113_/X vssd1 vssd1 vccd1 vccd1 _6323_/D sky130_fd_sc_hd__a31o_1
XFILLER_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6061_/B _6060_/B vssd1 vssd1 vccd1 vccd1 _6055_/A sky130_fd_sc_hd__nand2_1
X_3257_ _3257_/A vssd1 vssd1 vccd1 vccd1 _3257_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ input1/X vssd1 vssd1 vccd1 vccd1 _3313_/A sky130_fd_sc_hd__buf_2
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4821__B _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5829_ _5741_/A _5820_/A _5828_/X _5841_/B vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6053__C1 _5904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_452 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _5255_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__nand2_1
X_4091_ _4323_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ _5619_/A _5000_/B _4989_/A vssd1 vssd1 vccd1 vccd1 _4993_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3944_ _3944_/A _3944_/B vssd1 vssd1 vccd1 vccd1 _3972_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3875_ _3875_/A _3875_/B vssd1 vssd1 vccd1 vccd1 _3881_/B sky130_fd_sc_hd__xor2_1
X_5614_ _5614_/A _5622_/A vssd1 vssd1 vccd1 vccd1 _5616_/B sky130_fd_sc_hd__xnor2_1
X_6594_ _6594_/A _3314_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_5545_ _5575_/A _5575_/B _5543_/Y _5544_/X vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__a211o_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5476_ _5470_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5476_/X sky130_fd_sc_hd__and2b_1
X_4427_ _4427_/A _4427_/B vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__or2_1
XANTENNA__3273__A _3276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_A io_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4088__B _4088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4358_ _4358_/A _4358_/B vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__xnor2_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3309_ _3312_/A vssd1 vssd1 vccd1 vccd1 _3309_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4289_ _4297_/A _4297_/B _4288_/Y vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__a21bo_1
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6028_ _6299_/Q _6023_/X _6027_/X _6013_/X vssd1 vssd1 vccd1 vccd1 _6299_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_30 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5382__B _5382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4279__A _6281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4726__B _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _3659_/B _3659_/C _3659_/A vssd1 vssd1 vccd1 vccd1 _3664_/B sky130_fd_sc_hd__a21o_1
X_3591_ _3592_/A _3645_/C _3696_/B _4879_/B vssd1 vssd1 vccd1 vccd1 _3598_/B sky130_fd_sc_hd__a22o_1
X_5330_ _5330_/A _5485_/B _5330_/C vssd1 vssd1 vccd1 vccd1 _5370_/A sky130_fd_sc_hd__and3_1
XFILLER_55_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5261_ _5261_/A _5261_/B vssd1 vssd1 vccd1 vccd1 _5261_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4212_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4213_/B sky130_fd_sc_hd__or2_1
X_5192_ _5154_/B _5156_/X _5189_/Y _5546_/A vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__a211o_1
X_4143_ _4143_/A _4143_/B vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__xnor2_1
X_4074_ _5208_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4075_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4976_ _4961_/A _5000_/B _4961_/B _4974_/A vssd1 vssd1 vccd1 vccd1 _4977_/B sky130_fd_sc_hd__a22oi_1
X_3927_ _3928_/A _3928_/B _3928_/C vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3268__A _3270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3858_ _3903_/A vssd1 vssd1 vccd1 vccd1 _4960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3789_ _4929_/A _3947_/B vssd1 vssd1 vccd1 vccd1 _3885_/C sky130_fd_sc_hd__and2_1
X_6577_ _6577_/A _3288_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_5528_ _5621_/B _5629_/A _5621_/A vssd1 vssd1 vccd1 vccd1 _5622_/A sky130_fd_sc_hd__o21ai_1
XFILLER_105_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5459_ _5459_/A _5458_/A vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__or2b_1
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4546__B _4546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5219__A1_N _4059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4856_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _4832_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5287__B _5489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _4761_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__xor2_4
X_4692_ _4692_/A _4692_/B vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__nand2_1
X_3712_ _3668_/A _3668_/C _3668_/B vssd1 vssd1 vccd1 vccd1 _3713_/B sky130_fd_sc_hd__o21bai_1
X_6500_ _6500_/A _3204_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_3643_ _3643_/A _3643_/B vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__nand2_1
X_6362_ _6375_/CLK _6362_/D vssd1 vssd1 vccd1 vccd1 _6362_/Q sky130_fd_sc_hd__dfxtp_1
X_5313_ _5255_/A _5231_/D _5311_/X _5312_/X _5271_/X vssd1 vssd1 vccd1 vccd1 _5315_/A
+ sky130_fd_sc_hd__a32o_2
X_3574_ _3601_/A _3700_/B _3644_/B _4785_/A vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__a22o_1
XFILLER_114_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6293_ _6335_/CLK _6293_/D vssd1 vssd1 vccd1 vccd1 _6293_/Q sky130_fd_sc_hd__dfxtp_1
X_5244_ _5244_/A _5206_/X vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__or2b_1
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5175_ _5174_/A _5174_/B _5215_/A _5278_/B vssd1 vssd1 vccd1 vccd1 _5177_/B sky130_fd_sc_hd__a2bb2o_1
X_4126_ _4126_/A _4126_/B vssd1 vssd1 vccd1 vccd1 _4127_/B sky130_fd_sc_hd__xnor2_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4057_ _4009_/A _4008_/C _4008_/B vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _5183_/B vssd1 vssd1 vccd1 vccd1 _5000_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_7__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3290_ _3294_/A vssd1 vssd1 vccd1 vccd1 _3290_/Y sky130_fd_sc_hd__inv_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5931_ _5951_/A vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5862_ _5867_/A _5868_/A _5861_/X vssd1 vssd1 vccd1 vccd1 _5862_/Y sky130_fd_sc_hd__o21ai_1
X_4813_ _3645_/B _4879_/D _4787_/C _4707_/A vssd1 vssd1 vccd1 vccd1 _4818_/B sky130_fd_sc_hd__a22o_1
XFILLER_33_185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5793_ _5793_/A _5793_/B vssd1 vssd1 vccd1 vccd1 _5793_/X sky130_fd_sc_hd__or2_1
X_4744_ _4745_/B _4745_/C _4745_/A vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__o21a_1
X_4675_ _4877_/A _4877_/B _4675_/C _4785_/D vssd1 vssd1 vccd1 vccd1 _4712_/A sky130_fd_sc_hd__and4_1
X_3626_ _3626_/A _3626_/B vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__xor2_2
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6345_ _6345_/CLK _6345_/D vssd1 vssd1 vccd1 vccd1 _6345_/Q sky130_fd_sc_hd__dfxtp_1
X_3557_ _3483_/B _4814_/B _3400_/X _6286_/Q vssd1 vssd1 vccd1 vccd1 _3558_/B sky130_fd_sc_hd__o211a_1
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6276_ _6359_/CLK _6276_/D vssd1 vssd1 vccd1 vccd1 _6276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5227_ _5227_/A _5578_/A vssd1 vssd1 vccd1 vccd1 _5546_/C sky130_fd_sc_hd__nor2_1
X_3488_ _4651_/A _3600_/B _3643_/A _3487_/D vssd1 vssd1 vccd1 vccd1 _3489_/C sky130_fd_sc_hd__a22o_1
XANTENNA__3281__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5158_ _5158_/A _5158_/B vssd1 vssd1 vccd1 vccd1 _5159_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5089_ _5426_/B vssd1 vssd1 vccd1 vccd1 _5231_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4109_ _5165_/A _4365_/B _4365_/C vssd1 vssd1 vccd1 vccd1 _4114_/A sky130_fd_sc_hd__and3_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4788__A2 _4787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5001__A _5001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6162__A1 _5904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6561__77 vssd1 vssd1 vccd1 vccd1 _6561__77/HI _6561_/A sky130_fd_sc_hd__conb_1
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_496 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3191__A _3195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4460_ _4545_/A _4545_/B _4459_/Y vssd1 vssd1 vccd1 vccd1 _4593_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4391_ _4393_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _4392_/C sky130_fd_sc_hd__nor2_1
X_3411_ _3483_/B _4814_/B _3400_/X _6288_/Q vssd1 vssd1 vccd1 vccd1 _3548_/A sky130_fd_sc_hd__o211a_1
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3342_ _4731_/B vssd1 vssd1 vccd1 vccd1 _3505_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6130_ _6329_/Q _6146_/B vssd1 vssd1 vccd1 vccd1 _6131_/A sky130_fd_sc_hd__and2_1
XFILLER_112_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3276_/A vssd1 vssd1 vccd1 vccd1 _3273_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4197__A _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4561__A_N _4560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6061_ _6061_/A _6061_/B _6060_/B _6051_/A vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__or4bb_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5012_ _5012_/A _5032_/A vssd1 vssd1 vccd1 vccd1 _5013_/C sky130_fd_sc_hd__xor2_1
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5914_ _3333_/X _5896_/S _5912_/X _5913_/Y _6244_/A vssd1 vssd1 vccd1 vccd1 _5914_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5845_ _5690_/B _5757_/Y _5759_/X _5773_/B vssd1 vssd1 vccd1 vccd1 _5845_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5776_ _3333_/X _3384_/X _5775_/X vssd1 vssd1 vccd1 vccd1 _5776_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3276__A _3276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4727_ _4727_/A _4727_/B vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__nand2_2
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4658_ _4692_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__nand2_1
X_3609_ _4877_/D vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__clkbuf_2
X_4589_ _4589_/A _4595_/A vssd1 vssd1 vccd1 vccd1 _4589_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6328_ _6345_/CLK _6328_/D vssd1 vssd1 vccd1 vccd1 _6328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_466 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6259_ _6259_/A _6259_/B _6263_/C vssd1 vssd1 vccd1 vccd1 _6378_/D sky130_fd_sc_hd__nor3_1
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4697__A1 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5110__A2 _5145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3960_ _3960_/A _3960_/B vssd1 vssd1 vccd1 vccd1 _4010_/A sky130_fd_sc_hd__xor2_1
XANTENNA__4183__C _4337_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3891_ _3892_/A _3892_/B _3892_/C vssd1 vssd1 vccd1 vccd1 _3916_/A sky130_fd_sc_hd__o21ai_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5630_ _5630_/A _5630_/B vssd1 vssd1 vccd1 vccd1 _5634_/B sky130_fd_sc_hd__xnor2_1
X_5561_ _5561_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5683_/A sky130_fd_sc_hd__xnor2_2
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4512_ _4512_/A _4512_/B vssd1 vssd1 vccd1 vccd1 _4560_/A sky130_fd_sc_hd__xnor2_4
X_6525__44 vssd1 vssd1 vccd1 vccd1 _6525__44/HI _6525_/A sky130_fd_sc_hd__conb_1
X_5492_ _4266_/A _5365_/X _5468_/A _5491_/Y vssd1 vssd1 vccd1 vccd1 _5493_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4443_ _6274_/Q _4430_/B _4580_/B _5416_/A vssd1 vssd1 vccd1 vccd1 _4443_/X sky130_fd_sc_hd__a22o_1
X_4374_ _4374_/A _4374_/B vssd1 vssd1 vccd1 vccd1 _4378_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3325_ _5208_/A vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _6111_/X _6112_/X _6323_/Q _6201_/B vssd1 vssd1 vccd1 vccd1 _6113_/X sky130_fd_sc_hd__o211a_1
XFILLER_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3256_ _3257_/A vssd1 vssd1 vccd1 vccd1 _3256_/Y sky130_fd_sc_hd__inv_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6040_/A _6023_/X _6043_/X _6013_/X vssd1 vssd1 vccd1 vccd1 _6301_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_556 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5828_ _5690_/B _5793_/X _5792_/X _5773_/B vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5759_ _5759_/A _5759_/B vssd1 vssd1 vccd1 vccd1 _5759_/X sky130_fd_sc_hd__or2_1
XFILLER_108_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6300__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _5180_/C _3947_/B _4082_/B _4089_/Y vssd1 vssd1 vccd1 vccd1 _4098_/C sky130_fd_sc_hd__a31o_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4992_ _5023_/A _5024_/A vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__nand2_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3943_ _5129_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3819__A _3840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3874_ _3897_/A _3874_/B vssd1 vssd1 vccd1 vccd1 _3875_/B sky130_fd_sc_hd__and2_1
XFILLER_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5613_ _5613_/A _5613_/B vssd1 vssd1 vccd1 vccd1 _5618_/A sky130_fd_sc_hd__xnor2_1
X_6593_ _6593_/A _3312_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_5544_ _5308_/B _5544_/B vssd1 vssd1 vccd1 vccd1 _5544_/X sky130_fd_sc_hd__and2b_1
XFILLER_105_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5475_ _5483_/A _5483_/B vssd1 vssd1 vccd1 vccd1 _5478_/B sky130_fd_sc_hd__nand2_1
X_4426_ _4426_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4427_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4357_ _4463_/A _4463_/B vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__xor2_4
XFILLER_59_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4288_/A _4288_/B vssd1 vssd1 vccd1 vccd1 _4288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3308_ _3312_/A vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__inv_2
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3239_/A vssd1 vssd1 vccd1 vccd1 _3239_/Y sky130_fd_sc_hd__inv_2
X_6027_ _6027_/A _6027_/B _5989_/A vssd1 vssd1 vccd1 vccd1 _6027_/X sky130_fd_sc_hd__or3b_1
XFILLER_46_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6015__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3590_ _3580_/A _4898_/B _3589_/X vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__o21a_1
X_5260_ _5261_/A _5261_/B vssd1 vssd1 vccd1 vccd1 _5282_/B sky130_fd_sc_hd__xnor2_2
X_4211_ _5276_/A _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5191_ _5183_/C _5186_/B _5189_/Y _5190_/X vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__a211oi_2
X_4142_ _4142_/A _4142_/B _4142_/C vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__or3_1
X_4073_ _4365_/B _4365_/C vssd1 vssd1 vccd1 vccd1 _4396_/B sky130_fd_sc_hd__and2_2
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4933__A _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4975_ _4975_/A _4986_/A vssd1 vssd1 vccd1 vccd1 _4988_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3926_ _4484_/C _3924_/Y _3925_/X vssd1 vssd1 vccd1 vccd1 _3928_/C sky130_fd_sc_hd__o21a_1
XANTENNA__3549__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5467__C _5505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3857_ _5013_/A vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3788_ _5013_/A _4166_/B vssd1 vssd1 vccd1 vccd1 _3792_/A sky130_fd_sc_hd__nand2_1
X_6576_ _6576_/A _3286_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_5527_ _5527_/A _5527_/B vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3284__A _3288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5458_ _5458_/A _5459_/A vssd1 vssd1 vccd1 vccd1 _5462_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5389_ _5389_/A _5389_/B vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__xor2_2
X_4409_ _5484_/A _4409_/B _5484_/B vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__and3_1
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4282__A2 _4370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3194__A _3195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6567__83 vssd1 vssd1 vccd1 vccd1 _6567__83/HI _6567_/A sky130_fd_sc_hd__conb_1
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4760_ _4762_/A _4797_/A _4758_/A vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__a21o_2
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3711_ _3729_/A _3729_/B vssd1 vssd1 vccd1 vccd1 _3714_/B sky130_fd_sc_hd__xnor2_1
X_4691_ _4656_/Y _4659_/B _4657_/A vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__a21oi_1
XFILLER_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3642_ _3642_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__nand2_1
X_6361_ _6369_/CLK _6361_/D vssd1 vssd1 vccd1 vccd1 _6361_/Q sky130_fd_sc_hd__dfxtp_1
X_5312_ _5312_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__and3_1
X_3573_ _3696_/B vssd1 vssd1 vccd1 vccd1 _3644_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6292_ _6357_/CLK _6292_/D vssd1 vssd1 vccd1 vccd1 _6292_/Q sky130_fd_sc_hd__dfxtp_1
X_5243_ _5243_/A _5243_/B vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4928__A _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5174_ _5174_/A _5174_/B _4079_/A _5278_/B vssd1 vssd1 vccd1 vccd1 _5177_/A sky130_fd_sc_hd__or4bb_1
XANTENNA__3832__A _6278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4125_ _4117_/A _4117_/B _4145_/A vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__o21ai_1
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _4097_/A _4097_/B vssd1 vssd1 vccd1 vccd1 _4056_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3279__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4958_ _5038_/B vssd1 vssd1 vccd1 vccd1 _5183_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3909_ _4961_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _4484_/C sky130_fd_sc_hd__nand2_1
X_4889_ _4889_/A _4895_/A _4889_/C vssd1 vssd1 vccd1 vccd1 _4890_/C sky130_fd_sc_hd__nand3_1
XFILLER_20_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6559_ _6559_/A _3274_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4573__A _5001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3766__B2 _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4748__A _4787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5930_ _5951_/A vssd1 vssd1 vccd1 vccd1 _5930_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_120 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5861_ _6201_/B vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4812_ _4812_/A _4812_/B vssd1 vssd1 vccd1 vccd1 _4916_/B sky130_fd_sc_hd__xnor2_4
XFILLER_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5792_ _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__or2_1
X_4743_ _4743_/A _4743_/B vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__and2_1
X_4674_ _4645_/B _4675_/C _4785_/D _4645_/A vssd1 vssd1 vccd1 vccd1 _4674_/X sky130_fd_sc_hd__a22o_1
X_3625_ _3624_/A _3624_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3976_/C sky130_fd_sc_hd__a21o_1
X_6344_ _6345_/CLK _6344_/D vssd1 vssd1 vccd1 vccd1 _6344_/Q sky130_fd_sc_hd__dfxtp_1
X_3556_ _6288_/Q _3556_/B vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__nand2_4
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6275_ _6384_/CLK _6275_/D vssd1 vssd1 vccd1 vccd1 _6275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5226_ _5216_/X _5221_/B _5224_/A _5225_/X vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__o211a_1
X_3487_ _4664_/A _3600_/B _3643_/A _3487_/D vssd1 vssd1 vccd1 vccd1 _3643_/B sky130_fd_sc_hd__nand4_1
X_5157_ _5142_/A _5139_/B _5139_/C vssd1 vssd1 vccd1 vccd1 _5179_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4108_/A _4108_/B vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__or2_1
X_5088_ _5274_/C vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4039_ _4031_/A _4031_/B _4086_/A vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__a21o_1
XFILLER_16_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5001__B _5145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4568__A _5634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4390_ _5411_/A _4370_/B _4361_/C vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3410_ _3405_/X _3406_/X _6000_/A vssd1 vssd1 vccd1 vccd1 _4814_/B sky130_fd_sc_hd__a21oi_4
X_3341_ _4785_/A vssd1 vssd1 vccd1 vccd1 _4731_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5581__B _5672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3382__A _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3272_ _3276_/A vssd1 vssd1 vccd1 vccd1 _3272_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4197__B _4412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A _6060_/B _6060_/C vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__or3_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5011_ _5011_/A _5215_/B vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4925__B _5013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5913_ _5906_/A _5907_/X _5906_/B vssd1 vssd1 vccd1 vccd1 _5913_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5844_ _6380_/Q _5825_/Y _5835_/X _5838_/X _5843_/X vssd1 vssd1 vccd1 vccd1 _5844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5775_ _5769_/X _5684_/X _5771_/Y _4627_/Y _5774_/X vssd1 vssd1 vccd1 vccd1 _5775_/X
+ sky130_fd_sc_hd__a221o_1
X_4726_ _4726_/A _4726_/B _4726_/C vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__nand3_1
X_4657_ _4657_/A _4656_/Y vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__or2b_1
X_3608_ _4882_/A _3608_/B vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4588_ _4603_/B _4591_/B vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__nand2_1
X_6327_ _6345_/CLK _6327_/D vssd1 vssd1 vccd1 vccd1 _6327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_423 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3539_ _3551_/B vssd1 vssd1 vccd1 vccd1 _3762_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3292__A _3294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6258_ _6378_/Q _6258_/B _6258_/C vssd1 vssd1 vccd1 vccd1 _6263_/C sky130_fd_sc_hd__and3_1
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5209_ _5243_/A _5243_/B _5206_/X _5244_/A vssd1 vssd1 vccd1 vccd1 _5211_/B sky130_fd_sc_hd__a31o_1
X_6189_ _6351_/Q _6189_/B vssd1 vssd1 vccd1 vccd1 _6190_/A sky130_fd_sc_hd__and2_1
XFILLER_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4851__A _4865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_362 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3890_ _3890_/A _3905_/C vssd1 vssd1 vccd1 vccd1 _3892_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__5576__B _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__nor2_1
X_4511_ _5702_/A _4555_/A vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__and2b_1
X_5491_ _5491_/A vssd1 vssd1 vccd1 vccd1 _5491_/Y sky130_fd_sc_hd__clkinv_2
X_4442_ _5510_/A _4580_/B vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _4400_/A _4400_/B vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__or2_1
XFILLER_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3324_ _4194_/A vssd1 vssd1 vccd1 vccd1 _5208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6585__101 vssd1 vssd1 vccd1 vccd1 _6585__101/HI _6585_/A sky130_fd_sc_hd__conb_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6320_/Q _6319_/Q _6322_/Q _6321_/Q vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__or4_1
XFILLER_112_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3255_ _3257_/A vssd1 vssd1 vccd1 vccd1 _3255_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6043_/A _6043_/B _5989_/A vssd1 vssd1 vccd1 vccd1 _6043_/X sky130_fd_sc_hd__or3b_1
XANTENNA__3840__A _3840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_598 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5486__B _5486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3287__A _3288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5827_ _3383_/A _5826_/X _5820_/X _5733_/X vssd1 vssd1 vccd1 vccd1 _5827_/Y sky130_fd_sc_hd__a22oi_1
X_5758_ _5683_/B _5711_/B _5683_/A vssd1 vssd1 vccd1 vccd1 _5759_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4709_ _4877_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__nand2_1
X_5689_ _5779_/B _6302_/Q _5779_/A vssd1 vssd1 vccd1 vccd1 _5690_/B sky130_fd_sc_hd__or3b_2
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_410 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_58 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6053__A1 _6061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3197__A _3201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_62 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4731__D _4796_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3590__A2 _4898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6044__A1 _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4991_ _4983_/A _4991_/B vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__and2b_1
XFILLER_63_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3942_ _3973_/A vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3819__B _3840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3873_ _5037_/A _3950_/B _3906_/B _5001_/A vssd1 vssd1 vccd1 vccd1 _3874_/B sky130_fd_sc_hd__a22o_1
X_6592_ _6592_/A _3311_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_5612_ _5612_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5612_/X sky130_fd_sc_hd__or2_1
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5543_ _5578_/A _5578_/B _5578_/C vssd1 vssd1 vccd1 vccd1 _5543_/Y sky130_fd_sc_hd__nor3_1
X_5474_ _5474_/A vssd1 vssd1 vccd1 vccd1 _5483_/B sky130_fd_sc_hd__inv_2
XFILLER_105_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4425_ _4425_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__xor2_1
XANTENNA__6275__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4356_ _4356_/A _4356_/B vssd1 vssd1 vccd1 vccd1 _4463_/B sky130_fd_sc_hd__and2_2
XFILLER_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3307_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3312_/A sky130_fd_sc_hd__buf_8
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4288_/A _4288_/B vssd1 vssd1 vccd1 vccd1 _4297_/B sky130_fd_sc_hd__xor2_2
XFILLER_59_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6026_/A _6026_/B _6035_/B vssd1 vssd1 vccd1 vccd1 _6027_/B sky130_fd_sc_hd__and3_1
X_3238_ _3239_/A vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4576__A _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6298__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5573__C _5675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4210_ _5276_/A _4210_/B _4210_/C vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__and3_1
X_6510__29 vssd1 vssd1 vccd1 vccd1 _6510__29/HI _6510_/A sky130_fd_sc_hd__conb_1
XANTENNA__5870__A _5980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _5148_/X _5188_/X _5186_/A _5186_/Y vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__o211a_1
X_4141_ _4141_/A _4141_/B _4141_/C vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__and3_1
XFILLER_68_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4072_ _4072_/A _4072_/B _4072_/C vssd1 vssd1 vccd1 vccd1 _4365_/C sky130_fd_sc_hd__nand3_2
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4028__B1 _4367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4974_ _4974_/A _5000_/B vssd1 vssd1 vccd1 vccd1 _4986_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3925_ _4548_/A _4063_/B _3906_/B _4961_/A vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__a22o_1
X_3856_ _3793_/A _3793_/B _3855_/Y vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__a21o_1
X_6575_ _6575_/A _3287_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
X_3787_ _4131_/B vssd1 vssd1 vccd1 vccd1 _4166_/B sky130_fd_sc_hd__clkbuf_2
X_5526_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5527_/B sky130_fd_sc_hd__nor2_1
X_5457_ _5464_/A _5447_/B _5455_/X _5456_/X vssd1 vssd1 vccd1 vccd1 _5459_/A sky130_fd_sc_hd__a31oi_1
X_4408_ _4408_/A _4408_/B vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__xnor2_1
X_5388_ _5426_/A _5388_/B vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4339_ _4332_/A _4332_/B _4330_/X vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__o21a_1
XFILLER_115_78 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6009_ _6006_/X _6009_/B vssd1 vssd1 vccd1 vccd1 _6011_/A sky130_fd_sc_hd__and2b_1
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5955__A _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3475__A _3536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3710_ _3730_/B _3710_/B vssd1 vssd1 vccd1 vccd1 _3729_/B sky130_fd_sc_hd__nor2_1
X_4690_ _4663_/A _4662_/B _4689_/X vssd1 vssd1 vccd1 vccd1 _4701_/C sky130_fd_sc_hd__o21a_1
X_3641_ _3623_/A _3623_/B _3640_/X vssd1 vssd1 vccd1 vccd1 _3674_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__5584__B _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3572_ _3652_/B _3652_/C vssd1 vssd1 vccd1 vccd1 _3700_/B sky130_fd_sc_hd__and2_1
X_6582__98 vssd1 vssd1 vccd1 vccd1 _6582__98/HI _6582_/A sky130_fd_sc_hd__conb_1
X_6360_ _6369_/CLK _6360_/D vssd1 vssd1 vccd1 vccd1 _6360_/Q sky130_fd_sc_hd__dfxtp_1
X_5311_ _5312_/A _5444_/B _5444_/C _5246_/B _5274_/A vssd1 vssd1 vccd1 vccd1 _5311_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6291_ _6335_/CLK _6291_/D vssd1 vssd1 vccd1 vccd1 _6291_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _5242_/A _5242_/B vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__xor2_2
X_5173_ _5134_/A _5316_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5174_/B sky130_fd_sc_hd__a21oi_1
X_4124_ _4124_/A _4124_/B _4124_/C vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__or3_1
XFILLER_56_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4055_ _4055_/A _4055_/B vssd1 vssd1 vccd1 vccd1 _4097_/B sky130_fd_sc_hd__xor2_1
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4957_ _4966_/A _4957_/B vssd1 vssd1 vccd1 vccd1 _5038_/B sky130_fd_sc_hd__xnor2_4
X_3908_ _4925_/A vssd1 vssd1 vccd1 vccd1 _4961_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4888_ _4888_/A _4894_/A vssd1 vssd1 vccd1 vccd1 _4890_/B sky130_fd_sc_hd__or2b_1
XFILLER_32_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3839_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_552 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6558_ _6558_/A _3273_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5509_ _5621_/B _5509_/B vssd1 vssd1 vccd1 vccd1 _5628_/B sky130_fd_sc_hd__or2_1
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_20 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5685__A _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5860_ _6189_/B vssd1 vssd1 vccd1 vccd1 _6201_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4811_ _4918_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__xor2_4
XFILLER_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5791_ _6370_/Q _5791_/B vssd1 vssd1 vccd1 vccd1 _5791_/Y sky130_fd_sc_hd__nor2_1
X_4742_ _4742_/A _4742_/B vssd1 vssd1 vccd1 vccd1 _4743_/B sky130_fd_sc_hd__nand2_1
X_4673_ _4686_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4736_/A sky130_fd_sc_hd__xor2_1
X_3624_ _3624_/A _3624_/B _3624_/C vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__nand3_1
X_6343_ _6345_/CLK _6343_/D vssd1 vssd1 vccd1 vccd1 _6343_/Q sky130_fd_sc_hd__dfxtp_1
X_3555_ _3529_/B _3526_/C _3516_/Y vssd1 vssd1 vccd1 vccd1 _3560_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6274_ _6359_/CLK _6274_/D vssd1 vssd1 vccd1 vccd1 _6274_/Q sky130_fd_sc_hd__dfxtp_1
X_3486_ _4787_/A _3653_/B _3653_/C _3559_/B _6291_/Q vssd1 vssd1 vccd1 vccd1 _3487_/D
+ sky130_fd_sc_hd__a32o_1
X_5225_ _5186_/Y _5222_/X _5221_/A _5264_/A vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__a211o_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5156_ _5154_/A _5153_/C _5153_/B vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4107_ _4115_/A _4323_/B _4076_/C vssd1 vssd1 vccd1 vccd1 _4108_/B sky130_fd_sc_hd__a21oi_1
X_5087_ _5087_/A _5087_/B vssd1 vssd1 vccd1 vccd1 _5274_/C sky130_fd_sc_hd__xor2_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4038_ _4038_/A _4052_/B _4038_/C vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__and3_1
XANTENNA__5489__B _5489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3445__B2 _6291_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5989_ _5989_/A vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3753__A _5011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6552__68 vssd1 vssd1 vccd1 vccd1 _6552__68/HI _6552_/A sky130_fd_sc_hd__conb_1
X_3340_ _3592_/A vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__clkbuf_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__buf_6
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5010_ _5316_/B vssd1 vssd1 vccd1 vccd1 _5215_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5912_ _5906_/A _5901_/A _5907_/X _5899_/B vssd1 vssd1 vccd1 vccd1 _5912_/X sky130_fd_sc_hd__a31o_1
X_5843_ _5840_/Y _5842_/Y _5838_/X vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5774_ _5613_/A _5777_/B _5694_/X vssd1 vssd1 vccd1 vccd1 _5774_/X sky130_fd_sc_hd__a21o_1
X_4725_ _4726_/A _4726_/B _4726_/C vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__a21o_1
XFILLER_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4656_ _4656_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4656_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4155__A2 _4367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4587_ _4587_/A _4587_/B vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4669__A _4787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3607_ _3600_/Y _3632_/A _3602_/X vssd1 vssd1 vccd1 vccd1 _3608_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3538_ _3525_/Y _3534_/Y _3535_/Y _3536_/X vssd1 vssd1 vccd1 vccd1 _3543_/A sky130_fd_sc_hd__a211o_1
X_6326_ _6345_/CLK _6326_/D vssd1 vssd1 vccd1 vccd1 _6326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3469_ _3469_/A _3469_/B vssd1 vssd1 vccd1 vccd1 _3515_/B sky130_fd_sc_hd__xnor2_1
X_6257_ _6258_/B _6258_/C _6378_/Q vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__a21oi_1
X_5208_ _5208_/A _5246_/B _5251_/A vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__and3_1
X_6188_ _6188_/A vssd1 vssd1 vccd1 vccd1 _6351_/D sky130_fd_sc_hd__clkbuf_1
X_5139_ _5142_/A _5139_/B _5139_/C vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__nand3_1
XFILLER_69_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5812__C1 _6259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_444 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4510_ _4510_/A _4510_/B vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__xnor2_4
X_5490_ _5490_/A _5490_/B vssd1 vssd1 vccd1 vccd1 _5501_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5592__B _5637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4441_ _5936_/A _5349_/A _5450_/C vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__and3_2
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4372_ _4372_/A _4372_/B vssd1 vssd1 vccd1 vccd1 _4400_/B sky130_fd_sc_hd__xor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6316_/Q _6315_/Q _6318_/Q _6317_/Q vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__or4_1
XFILLER_112_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3323_ _5328_/A vssd1 vssd1 vccd1 vccd1 _4194_/A sky130_fd_sc_hd__clkbuf_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3257_/A vssd1 vssd1 vccd1 vccd1 _3254_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6042_/A _6042_/B _6042_/C vssd1 vssd1 vccd1 vccd1 _6043_/B sky130_fd_sc_hd__and3_1
XANTENNA__3840__B _3840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5826_ _5813_/X _5724_/Y _5727_/Y _5814_/X vssd1 vssd1 vccd1 vccd1 _5826_/X sky130_fd_sc_hd__a22o_1
X_5757_ _5757_/A _5757_/B vssd1 vssd1 vccd1 vccd1 _5757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4708_ _4842_/B _4707_/X _4719_/A vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__a21boi_1
X_6516__35 vssd1 vssd1 vccd1 vccd1 _6516__35/HI _6516_/A sky130_fd_sc_hd__conb_1
XFILLER_108_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5688_ _5779_/A _5701_/B _6302_/Q vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__or3b_2
X_4639_ _4768_/C vssd1 vssd1 vccd1 vccd1 _4675_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6309_ _6384_/CLK _6309_/D vssd1 vssd1 vccd1 vccd1 _6309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4064__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4990_ _5023_/B _5024_/A vssd1 vssd1 vccd1 vccd1 _4997_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5587__B _5637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3941_ _3941_/A _3975_/A vssd1 vssd1 vccd1 vccd1 _3973_/A sky130_fd_sc_hd__xor2_1
X_3872_ _5059_/A vssd1 vssd1 vccd1 vccd1 _5001_/A sky130_fd_sc_hd__buf_2
XFILLER_90_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6591_ _6591_/A _3310_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_5611_ _5664_/A _5664_/B _5610_/X vssd1 vssd1 vccd1 vccd1 _5612_/B sky130_fd_sc_hd__o21a_1
X_5542_ _5582_/A _5582_/B _5541_/X vssd1 vssd1 vccd1 vccd1 _5575_/B sky130_fd_sc_hd__a21o_2
X_5473_ _5473_/A _5473_/B vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__xnor2_1
X_4424_ _4455_/A _4455_/B _4423_/X vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__o21ai_1
X_4355_ _4358_/A _4358_/B vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__or2b_1
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _3306_/A vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4286_ _4309_/A _4309_/B _4285_/A vssd1 vssd1 vccd1 vccd1 _4288_/B sky130_fd_sc_hd__o21bai_2
XFILLER_58_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3239_/A vssd1 vssd1 vccd1 vccd1 _3237_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6026_/A _6026_/B _6035_/B vssd1 vssd1 vccd1 vccd1 _6027_/A sky130_fd_sc_hd__a21oi_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3298__A _3300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5809_ _6372_/Q _5805_/B _5808_/X _6373_/Q vssd1 vssd1 vccd1 vccd1 _5809_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _4142_/A _4142_/B _4142_/C vssd1 vssd1 vccd1 vccd1 _4141_/C sky130_fd_sc_hd__o21ai_4
XFILLER_68_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _4365_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4973_ _5003_/A _5003_/B vssd1 vssd1 vccd1 vccd1 _4998_/B sky130_fd_sc_hd__and2_1
XFILLER_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5776__A1 _3333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3924_ _4548_/A _4484_/B vssd1 vssd1 vccd1 vccd1 _3924_/Y sky130_fd_sc_hd__nand2_1
X_3855_ _3939_/A _3939_/B vssd1 vssd1 vccd1 vccd1 _3855_/Y sky130_fd_sc_hd__nor2_1
X_3786_ _3786_/A vssd1 vssd1 vccd1 vccd1 _4131_/B sky130_fd_sc_hd__clkbuf_2
X_6574_ _6574_/A _3290_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_5525_ _5628_/B _5525_/B vssd1 vssd1 vccd1 vccd1 _5629_/A sky130_fd_sc_hd__and2b_1
X_5456_ _5454_/A _5456_/B vssd1 vssd1 vccd1 vccd1 _5456_/X sky130_fd_sc_hd__and2b_1
X_4407_ _4459_/A _4459_/B vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__xor2_1
X_5387_ _5404_/C _5387_/B vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__xnor2_2
XFILLER_115_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4338_/A _4352_/B vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__xor2_1
XANTENNA__4396__B _4396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A io_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4269_ _5386_/A _4324_/B _4268_/C vssd1 vssd1 vccd1 vccd1 _4270_/B sky130_fd_sc_hd__a21oi_1
X_6008_ _6297_/Q _6031_/B vssd1 vssd1 vccd1 vccd1 _6009_/B sky130_fd_sc_hd__or2_1
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3475__B _3536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3545_/B _3640_/B vssd1 vssd1 vccd1 vccd1 _3640_/X sky130_fd_sc_hd__and2b_1
X_3571_ _4879_/B vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__buf_2
X_5310_ _5310_/A _5310_/B vssd1 vssd1 vccd1 vccd1 _5541_/B sky130_fd_sc_hd__xnor2_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6290_ _6335_/CLK _6290_/D vssd1 vssd1 vccd1 vccd1 _6290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5241_ _5281_/A _5281_/B vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__and2_1
XFILLER_102_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5172_ _5195_/A _5172_/B _5172_/C vssd1 vssd1 vccd1 vccd1 _5174_/A sky130_fd_sc_hd__and3_2
X_4123_ _5199_/A _4210_/B _4122_/C _4122_/D vssd1 vssd1 vccd1 vccd1 _4124_/C sky130_fd_sc_hd__a22oi_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4054_ _4063_/C _4054_/B vssd1 vssd1 vccd1 vccd1 _4055_/B sky130_fd_sc_hd__xnor2_2
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4956_ _4941_/Y _4944_/B _4942_/A vssd1 vssd1 vccd1 vccd1 _4957_/B sky130_fd_sc_hd__a21o_1
X_6558__74 vssd1 vssd1 vccd1 vccd1 _6558__74/HI _6558_/A sky130_fd_sc_hd__conb_1
X_3907_ _4974_/A _4138_/B vssd1 vssd1 vccd1 vccd1 _3922_/A sky130_fd_sc_hd__nand2_1
X_4887_ _4889_/A _4889_/C _4895_/A vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__a21o_1
X_3838_ _5133_/A vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6557_ _6557_/A _3272_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
X_3769_ _3810_/B _3769_/B vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__nand2_1
X_5508_ _5508_/A _5508_/B vssd1 vssd1 vccd1 vccd1 _5509_/B sky130_fd_sc_hd__and2_1
XFILLER_105_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5439_ _6277_/Q _5439_/B vssd1 vssd1 vccd1 vccd1 _5440_/C sky130_fd_sc_hd__and2_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_190 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6288__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5031__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5966__A _5966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5912__A1 _5906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4810_ _4810_/A _4810_/B vssd1 vssd1 vccd1 vccd1 _4918_/B sky130_fd_sc_hd__and2_2
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5790_ _6241_/B _5787_/B _5791_/B _6370_/Q vssd1 vssd1 vccd1 vccd1 _5790_/Y sky130_fd_sc_hd__a22oi_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4747_/B _4747_/A vssd1 vssd1 vccd1 vccd1 _4745_/C sky130_fd_sc_hd__and2b_1
X_4672_ _5955_/A _4726_/B vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__nand2_1
X_3623_ _3623_/A _3623_/B vssd1 vssd1 vccd1 vccd1 _3941_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4706__A2 _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6342_ _6345_/CLK _6342_/D vssd1 vssd1 vccd1 vccd1 _6342_/Q sky130_fd_sc_hd__dfxtp_1
X_3554_ _3552_/A _3575_/C _3553_/Y vssd1 vssd1 vccd1 vccd1 _3570_/A sky130_fd_sc_hd__a21o_1
XFILLER_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6273_ _6383_/Q _6270_/B _6272_/Y vssd1 vssd1 vccd1 vccd1 _6383_/D sky130_fd_sc_hd__o21a_1
X_3485_ _3516_/A vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5224_ _5224_/A vssd1 vssd1 vccd1 vccd1 _5227_/A sky130_fd_sc_hd__inv_2
XFILLER_111_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6491__10 vssd1 vssd1 vccd1 vccd1 _6491__10/HI _6491_/A sky130_fd_sc_hd__conb_1
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _5550_/A _5550_/B _5550_/C vssd1 vssd1 vccd1 vccd1 _5596_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4106_ _4106_/A _4106_/B vssd1 vssd1 vccd1 vccd1 _4139_/B sky130_fd_sc_hd__xnor2_1
X_5086_ _5086_/A _5086_/B vssd1 vssd1 vccd1 vccd1 _5103_/A sky130_fd_sc_hd__xnor2_1
X_4037_ _4079_/A _3786_/A _4052_/A _4036_/D vssd1 vssd1 vccd1 vccd1 _4038_/C sky130_fd_sc_hd__a22o_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5988_ _6023_/A vssd1 vssd1 vccd1 vccd1 _5988_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4939_ _4954_/A _4939_/B vssd1 vssd1 vccd1 vccd1 _4941_/B sky130_fd_sc_hd__and2_1
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3753__B _4168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4865__A _4865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6303__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3270_ _3270_/A vssd1 vssd1 vccd1 vccd1 _3270_/Y sky130_fd_sc_hd__inv_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5911_ _5906_/A _5857_/X _5910_/Y _5872_/X vssd1 vssd1 vccd1 vccd1 _6280_/D sky130_fd_sc_hd__o211a_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5842_ _5841_/Y _5837_/Y _6379_/Q vssd1 vssd1 vccd1 vccd1 _5842_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5773_ _5773_/A _5773_/B vssd1 vssd1 vccd1 vccd1 _5777_/B sky130_fd_sc_hd__nand2_1
X_4724_ _4718_/A _4718_/B _4715_/X vssd1 vssd1 vccd1 vccd1 _4726_/C sky130_fd_sc_hd__o21a_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4655_ _4656_/A _4654_/X _4656_/B vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__a21oi_1
X_4586_ _5646_/A _4586_/B vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__xor2_1
X_3606_ _3629_/B _3606_/B vssd1 vssd1 vccd1 vccd1 _3634_/B sky130_fd_sc_hd__or2_1
X_3537_ _3525_/Y _3534_/Y _3535_/Y _3536_/X vssd1 vssd1 vccd1 vccd1 _3544_/A sky130_fd_sc_hd__a211oi_1
X_6325_ _6345_/CLK _6325_/D vssd1 vssd1 vccd1 vccd1 _6325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_114 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6256_ _6258_/B _6258_/C _6255_/Y vssd1 vssd1 vccd1 vccd1 _6377_/D sky130_fd_sc_hd__o21a_1
X_3468_ _3516_/A _3522_/B _4818_/A vssd1 vssd1 vccd1 vccd1 _3514_/B sky130_fd_sc_hd__a21boi_1
X_5207_ _5294_/A _5469_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5251_/A sky130_fd_sc_hd__and3_1
X_3399_ _6298_/Q _3449_/A _3401_/A vssd1 vssd1 vccd1 vccd1 _3549_/B sky130_fd_sc_hd__or3_1
X_6187_ _6187_/A input6/X vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__and2_1
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5138_ _5138_/A _5138_/B vssd1 vssd1 vccd1 vccd1 _5139_/C sky130_fd_sc_hd__xor2_1
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5069_ _5070_/A _5070_/B vssd1 vssd1 vccd1 vccd1 _5071_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4579__B _5511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6140__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4440_ _4440_/A _4440_/B vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__xnor2_1
X_4371_ _5382_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4372_/B sky130_fd_sc_hd__nand2_1
X_6110_ _6316_/Q _6317_/Q _6110_/C vssd1 vssd1 vccd1 vccd1 _6110_/X sky130_fd_sc_hd__and3_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3322_ _6281_/Q vssd1 vssd1 vccd1 vccd1 _5328_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3253_ _3257_/A vssd1 vssd1 vccd1 vccd1 _3253_/Y sky130_fd_sc_hd__inv_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6042_/A _6042_/B _6042_/C vssd1 vssd1 vccd1 vccd1 _6043_/A sky130_fd_sc_hd__a21oi_1
XFILLER_112_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5825_ _5890_/A _5820_/X _5824_/X _3384_/X vssd1 vssd1 vccd1 vccd1 _5825_/Y sky130_fd_sc_hd__a22oi_2
X_5756_ _5710_/A _5710_/B _4626_/A vssd1 vssd1 vccd1 vccd1 _5757_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4707_ _4707_/A _4707_/B _4768_/D vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__and3_1
X_5687_ _6061_/A _5770_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _5687_/X sky130_fd_sc_hd__o21a_1
X_4638_ _4638_/A _4638_/B vssd1 vssd1 vccd1 vccd1 _4680_/A sky130_fd_sc_hd__or2_1
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4569_ _4569_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6308_ _6369_/CLK _6308_/D vssd1 vssd1 vccd1 vccd1 _6308_/Q sky130_fd_sc_hd__dfxtp_1
X_6239_ _6242_/A _6239_/B vssd1 vssd1 vccd1 vccd1 _6239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3940_ _5091_/A _3940_/B vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__nand2_1
XFILLER_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6045__A _6061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3871_ _4088_/B vssd1 vssd1 vccd1 vccd1 _3950_/B sky130_fd_sc_hd__clkbuf_2
X_6590_ _6590_/A _3309_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5610_ _5676_/A _5610_/B vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__or2_1
X_5541_ _5346_/B _5541_/B vssd1 vssd1 vccd1 vccd1 _5541_/X sky130_fd_sc_hd__and2b_1
X_5472_ _5472_/A _5472_/B vssd1 vssd1 vccd1 vccd1 _5483_/A sky130_fd_sc_hd__xor2_1
X_4423_ _4423_/A _4423_/B vssd1 vssd1 vccd1 vccd1 _4423_/X sky130_fd_sc_hd__or2_1
X_4354_ _4354_/A _4354_/B vssd1 vssd1 vccd1 vccd1 _4358_/B sky130_fd_sc_hd__xnor2_1
X_3305_ _3306_/A vssd1 vssd1 vccd1 vccd1 _3305_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4285_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4309_/B sky130_fd_sc_hd__or2_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _6299_/Q _6031_/B vssd1 vssd1 vccd1 vccd1 _6035_/B sky130_fd_sc_hd__xor2_1
X_3236_ _3239_/A vssd1 vssd1 vccd1 vccd1 _3236_/Y sky130_fd_sc_hd__inv_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5808_ _5755_/A _5778_/X _5807_/X _5706_/X vssd1 vssd1 vccd1 vccd1 _5808_/X sky130_fd_sc_hd__o2bb2a_1
X_5739_ _5736_/X _5738_/X _5777_/A vssd1 vssd1 vccd1 vccd1 _5739_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_592 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5846__A1_N _5755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__xor2_1
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A _4972_/B vssd1 vssd1 vccd1 vccd1 _5003_/B sky130_fd_sc_hd__xnor2_1
XFILLER_63_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _4978_/A _4484_/B _3923_/C vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__and3_1
X_3854_ _3854_/A _3879_/C vssd1 vssd1 vccd1 vccd1 _3939_/B sky130_fd_sc_hd__xor2_1
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3785_ _3840_/A _3785_/B vssd1 vssd1 vccd1 vccd1 _3786_/A sky130_fd_sc_hd__nand2_1
X_6573_ _6573_/A _3292_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_5524_ _5642_/A _5635_/B _5523_/A vssd1 vssd1 vccd1 vccd1 _5525_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4958__A _5038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5455_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5455_/X sky130_fd_sc_hd__or2_1
X_4406_ _4408_/A _4408_/B _4405_/Y vssd1 vssd1 vccd1 vccd1 _4459_/B sky130_fd_sc_hd__a21oi_1
X_5386_ _5386_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__nand2_1
X_4337_ _5489_/A _4337_/B _4337_/C vssd1 vssd1 vccd1 vccd1 _4352_/B sky130_fd_sc_hd__and3_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _5386_/A _4268_/B _4268_/C vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__and3_1
XFILLER_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3219_ _3220_/A vssd1 vssd1 vccd1 vccd1 _3219_/Y sky130_fd_sc_hd__inv_2
X_6007_ _6016_/B vssd1 vssd1 vccd1 vccd1 _6031_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4199_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__or2_1
XFILLER_39_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5699__A _5819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3947__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3570_/A _3570_/B vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__xnor2_2
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5143__B1 _4062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5240_ _5264_/A _5264_/B vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__nor2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5171_ _5230_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5172_/C sky130_fd_sc_hd__and2_1
XFILLER_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4122_ _5255_/A _4122_/B _4122_/C _4122_/D vssd1 vssd1 vccd1 vccd1 _4124_/B sky130_fd_sc_hd__and4_1
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4053_ _4053_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _4054_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_4__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4955_ _4954_/A _4953_/B _4954_/Y vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__o21ai_4
XFILLER_52_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3906_ _4960_/A _3906_/B vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__nand2_1
X_4886_ _4894_/A _4894_/B _4894_/C vssd1 vssd1 vccd1 vccd1 _4895_/A sky130_fd_sc_hd__a21oi_2
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3837_ _5230_/A vssd1 vssd1 vccd1 vccd1 _5133_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6556_ _6556_/A _3270_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
X_3768_ _3768_/A _3768_/B vssd1 vssd1 vccd1 vccd1 _3769_/B sky130_fd_sc_hd__nand2_1
X_6573__89 vssd1 vssd1 vccd1 vccd1 _6573__89/HI _6573_/A sky130_fd_sc_hd__conb_1
X_5507_ _5508_/A _5508_/B vssd1 vssd1 vccd1 vccd1 _5621_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3699_ _4877_/A _3503_/A _3503_/B _3644_/B _4796_/A vssd1 vssd1 vccd1 vccd1 _3700_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_105_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5438_ _5484_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5452_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5369_ _5369_/A _5369_/B vssd1 vssd1 vccd1 vccd1 _5390_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5031__B _5358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5912__A2 _5901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4732_/A _4755_/A _4727_/A vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__o21ai_4
XFILLER_14_381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4671_ _4677_/A _4677_/B _4666_/X vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__3396__B _6060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3622_ _3624_/B _3624_/C _3624_/A vssd1 vssd1 vccd1 vccd1 _3623_/B sky130_fd_sc_hd__a21bo_1
X_6341_ _6345_/CLK _6341_/D vssd1 vssd1 vccd1 vccd1 _6341_/Q sky130_fd_sc_hd__dfxtp_1
X_3553_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3553_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6272_ _6383_/Q _6270_/B _6218_/A vssd1 vssd1 vccd1 vccd1 _6272_/Y sky130_fd_sc_hd__a21oi_1
X_3484_ _3484_/A _3580_/A _3653_/C _3458_/A vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__or4bb_1
XFILLER_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5223_ _5221_/A _5264_/A _5186_/Y _5222_/X vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__o211ai_2
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5550_/C sky130_fd_sc_hd__nand2_1
X_4105_ _4105_/A _4105_/B vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5419__A1 _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _5085_/A _5215_/B vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4036_ _5215_/A _4131_/B _4052_/A _4036_/D vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__nand4_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4971__A _5634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5987_ _5989_/A vssd1 vssd1 vccd1 vccd1 _6023_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4938_ _4937_/A _4937_/B _4936_/X vssd1 vssd1 vccd1 vccd1 _4939_/B sky130_fd_sc_hd__o21bai_1
X_4869_ _4869_/A _4869_/B _4869_/C vssd1 vssd1 vccd1 vccd1 _4889_/A sky130_fd_sc_hd__nand3_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6539_ _6539_/A _3250_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5910_ _5910_/A _5910_/B vssd1 vssd1 vccd1 vccd1 _5910_/Y sky130_fd_sc_hd__nand2_1
X_5841_ _5885_/A _5841_/B vssd1 vssd1 vccd1 vccd1 _5841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5772_ _5813_/B _5779_/B _5814_/C vssd1 vssd1 vccd1 vccd1 _5773_/B sky130_fd_sc_hd__or3b_2
XANTENNA__3200__A _3201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4723_ _4733_/B _4733_/C _4733_/A vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4654_ _4644_/A _4693_/A _4692_/B _4694_/A vssd1 vssd1 vccd1 vccd1 _4654_/X sky130_fd_sc_hd__a22o_1
X_6543__59 vssd1 vssd1 vccd1 vccd1 _6543__59/HI _6543_/A sky130_fd_sc_hd__conb_1
X_4585_ _5001_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4585_/Y sky130_fd_sc_hd__xnor2_1
X_3605_ _3604_/B _3605_/B vssd1 vssd1 vccd1 vccd1 _3606_/B sky130_fd_sc_hd__and2b_1
X_3536_ _3536_/A _3536_/B _3536_/C vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__and3_1
X_6324_ _6345_/CLK _6324_/D vssd1 vssd1 vccd1 vccd1 _6324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6255_ _6258_/B _6258_/C _6218_/A vssd1 vssd1 vccd1 vccd1 _6255_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5206_ _5208_/A _5489_/B _5166_/C vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3467_ _6290_/Q _3556_/B vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__nand2_2
X_6186_ _6343_/Q _6344_/Q _5861_/X _6182_/X _6185_/X vssd1 vssd1 vccd1 vccd1 _6350_/D
+ sky130_fd_sc_hd__a41o_1
X_3398_ _6304_/Q _6303_/Q _6297_/Q vssd1 vssd1 vccd1 vccd1 _3401_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5137_ _5136_/A _5136_/B _5180_/C _5236_/B vssd1 vssd1 vccd1 vccd1 _5139_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _5129_/A _5388_/B vssd1 vssd1 vccd1 vccd1 _5070_/B sky130_fd_sc_hd__nand2_2
X_4019_ _4019_/A vssd1 vssd1 vccd1 vccd1 _4271_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6140__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4370_ _5246_/A _4370_/B vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__nand2_1
X_3321_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3321_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3252_ _3258_/A vssd1 vssd1 vccd1 vccd1 _3257_/A sky130_fd_sc_hd__buf_8
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6046_/B vssd1 vssd1 vccd1 vccd1 _6042_/C sky130_fd_sc_hd__xor2_1
XFILLER_79_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5824_ _5813_/X _5710_/X _5711_/Y _5814_/X vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__a22o_1
X_6592__108 vssd1 vssd1 vccd1 vccd1 _6592__108/HI _6592_/A sky130_fd_sc_hd__conb_1
X_5755_ _5755_/A vssd1 vssd1 vccd1 vccd1 _5901_/A sky130_fd_sc_hd__clkbuf_2
X_5686_ _5779_/B vssd1 vssd1 vccd1 vccd1 _6061_/A sky130_fd_sc_hd__clkbuf_2
X_4706_ _3592_/A _4707_/B _4641_/A _3522_/A vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__a22o_1
X_4637_ _4846_/B _4694_/A _3484_/A _4814_/C vssd1 vssd1 vccd1 vccd1 _4638_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_116_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4568_ _5634_/A vssd1 vssd1 vccd1 vccd1 _5899_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4499_ _4487_/A _4499_/B _4499_/C _4499_/D vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__and4b_2
X_6307_ _6384_/CLK _6307_/D vssd1 vssd1 vccd1 vccd1 _6307_/Q sky130_fd_sc_hd__dfxtp_1
X_3519_ _3386_/A _3391_/A _5993_/A vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__a21oi_4
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6238_ _6241_/B _6241_/C vssd1 vssd1 vccd1 vccd1 _6239_/B sky130_fd_sc_hd__and2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6344_/D sky130_fd_sc_hd__clkbuf_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6507__26 vssd1 vssd1 vccd1 vccd1 _6507__26/HI _6507_/A sky130_fd_sc_hd__conb_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3870_ _3870_/A _3901_/A vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__or2_1
XFILLER_16_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5540_ _5586_/A _5586_/B _5539_/X vssd1 vssd1 vccd1 vccd1 _5582_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6061__A _6061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5471_ _5471_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5472_/B sky130_fd_sc_hd__and3_1
X_4422_ _4423_/A _4423_/B vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__xnor2_1
X_6521__40 vssd1 vssd1 vccd1 vccd1 _6521__40/HI _6521_/A sky130_fd_sc_hd__conb_1
XFILLER_98_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4353_ _4353_/A _4353_/B vssd1 vssd1 vccd1 vccd1 _4358_/A sky130_fd_sc_hd__nor2_1
X_3304_ _3306_/A vssd1 vssd1 vccd1 vccd1 _3304_/Y sky130_fd_sc_hd__inv_2
X_4284_ _4283_/B _4284_/B vssd1 vssd1 vccd1 vccd1 _4285_/B sky130_fd_sc_hd__and2b_1
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _3239_/A vssd1 vssd1 vccd1 vccd1 _3235_/Y sky130_fd_sc_hd__inv_2
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _6023_/A vssd1 vssd1 vccd1 vccd1 _6023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3999_ _5314_/A vssd1 vssd1 vccd1 vccd1 _5276_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5807_ _5690_/A _5759_/X _5815_/B _5757_/Y vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4754__B2 _5325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3557__A2 _4814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5738_ _5815_/A _5792_/A _5792_/B vssd1 vssd1 vccd1 vccd1 _5738_/X sky130_fd_sc_hd__or3_1
XFILLER_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5669_ _5669_/A _5669_/B vssd1 vssd1 vccd1 vccd1 _5669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6579__95 vssd1 vssd1 vccd1 vccd1 _6579__95/HI _6579_/A sky130_fd_sc_hd__conb_1
XANTENNA__4993__A1 _5619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4113__B _4340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5170__A1 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _5634_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__and2_1
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3922_ _3922_/A _4484_/C vssd1 vssd1 vccd1 vccd1 _3928_/A sky130_fd_sc_hd__nor2_1
X_3853_ _3961_/B _3870_/A vssd1 vssd1 vccd1 vccd1 _3879_/C sky130_fd_sc_hd__xor2_1
XFILLER_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3784_ _3782_/A _3782_/B _3781_/X vssd1 vssd1 vccd1 vccd1 _3785_/B sky130_fd_sc_hd__o21bai_2
X_6572_ _6572_/A _3294_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_5523_ _5523_/A _5523_/B vssd1 vssd1 vccd1 vccd1 _5635_/B sky130_fd_sc_hd__nand2_1
X_6498__17 vssd1 vssd1 vccd1 vccd1 _6498__17/HI _6498_/A sky130_fd_sc_hd__conb_1
X_5454_ _5454_/A _5456_/B vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5385_ _5383_/A _5383_/B _5384_/X vssd1 vssd1 vccd1 vccd1 _5404_/C sky130_fd_sc_hd__a21o_1
X_4405_ _4405_/A _4405_/B vssd1 vssd1 vccd1 vccd1 _4405_/Y sky130_fd_sc_hd__nor2_1
X_4336_ _4353_/A _4336_/B vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__or2_1
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _4227_/B _4303_/A _4274_/A _4274_/B vssd1 vssd1 vccd1 vccd1 _4268_/C sky130_fd_sc_hd__o22ai_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3218_ _3220_/A vssd1 vssd1 vccd1 vccd1 _3218_/Y sky130_fd_sc_hd__inv_2
X_4198_ _4198_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6006_ _6297_/Q _6016_/B vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__and2_1
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3947__B _3947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5915__B1 _3333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5170_ _5085_/A _5404_/B _5202_/B _5169_/A vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__a31o_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4121_ _5195_/A _3940_/B _4120_/X vssd1 vssd1 vccd1 vccd1 _4122_/D sky130_fd_sc_hd__a21o_1
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4052_ _4052_/A _4052_/B vssd1 vssd1 vccd1 vccd1 _4063_/C sky130_fd_sc_hd__nand2_1
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3457__A1 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4954_ _4954_/A _4954_/B vssd1 vssd1 vccd1 vccd1 _4954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3905_ _4978_/A _4063_/B _3905_/C vssd1 vssd1 vccd1 vccd1 _3913_/B sky130_fd_sc_hd__and3_1
X_4885_ _4885_/A _4885_/B vssd1 vssd1 vccd1 vccd1 _4894_/C sky130_fd_sc_hd__or2_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3836_ _5231_/A vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4969__A _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3767_ _3768_/A _3768_/B vssd1 vssd1 vccd1 vccd1 _3810_/B sky130_fd_sc_hd__or2_1
X_6555_ _6555_/A _3269_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_5506_ _5519_/B _5520_/B _5519_/A vssd1 vssd1 vccd1 vccd1 _5508_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__3592__B _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3698_ _4787_/A vssd1 vssd1 vccd1 vccd1 _4877_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5437_ _5437_/A vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__inv_2
XFILLER_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5368_ _5246_/A _5365_/X _5392_/B _5367_/X vssd1 vssd1 vccd1 vccd1 _5369_/B sky130_fd_sc_hd__a31o_1
X_5299_ _5318_/A _5318_/B _5298_/A vssd1 vssd1 vccd1 vccd1 _5302_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4319_ _4320_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__xor2_1
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5312__B _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6549__65 vssd1 vssd1 vccd1 vccd1 _6549__65/HI _6549_/A sky130_fd_sc_hd__conb_1
XFILLER_23_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4731_/A _4864_/C vssd1 vssd1 vccd1 vccd1 _4677_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3621_ _3621_/A _3621_/B _3621_/C vssd1 vssd1 vccd1 vccd1 _3624_/A sky130_fd_sc_hd__or3_1
XANTENNA__3693__A _3693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6340_ _6357_/CLK _6340_/D vssd1 vssd1 vccd1 vccd1 _6340_/Q sky130_fd_sc_hd__dfxtp_1
X_3552_ _3552_/A _3575_/C vssd1 vssd1 vccd1 vccd1 _3562_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6271_ _6382_/Q _6267_/B _6270_/Y vssd1 vssd1 vccd1 vccd1 _6382_/D sky130_fd_sc_hd__o21a_1
X_3483_ _4814_/A _3483_/B _3436_/B vssd1 vssd1 vccd1 vccd1 _3580_/A sky130_fd_sc_hd__or3b_2
XFILLER_102_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5186_/B _5186_/C _5186_/D _5186_/A vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5153_ _5154_/A _5153_/B _5153_/C vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__nand3_1
XFILLER_69_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4104_ _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__xor2_4
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_408 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5084_ _5075_/A _5075_/B _5075_/C vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4627__B1 _4516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4035_ _5133_/A _4210_/B _3987_/B _5134_/A vssd1 vssd1 vccd1 vccd1 _4036_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3868__A _4051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6244__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5986_ _5982_/X _5983_/Y _5984_/X _5985_/X vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__o22a_1
X_4937_ _4937_/A _4937_/B _4936_/X vssd1 vssd1 vccd1 vccd1 _4954_/A sky130_fd_sc_hd__or3b_2
X_4868_ _4868_/A _4868_/B _4868_/C vssd1 vssd1 vccd1 vccd1 _4869_/C sky130_fd_sc_hd__nand3_1
XFILLER_20_330 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3819_ _3840_/A _3840_/B vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__nor2_2
X_4799_ _4818_/A _4800_/B vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__and2_1
XFILLER_21_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6538_ _6538_/A _3249_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_21_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5034__B1 _5355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6064__A _6254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5840_ _3384_/A _5826_/X _5820_/X _5733_/X _5839_/Y vssd1 vssd1 vccd1 vccd1 _5840_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_15_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ _6063_/A _6061_/A _6061_/B vssd1 vssd1 vccd1 vccd1 _5771_/Y sky130_fd_sc_hd__nor3_2
X_4722_ _4722_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__xor2_1
XFILLER_21_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4653_ _5966_/A _4694_/C _4693_/A vssd1 vssd1 vccd1 vccd1 _4656_/A sky130_fd_sc_hd__or3b_1
X_4584_ _5646_/A _4586_/B _4583_/Y vssd1 vssd1 vccd1 vccd1 _4584_/Y sky130_fd_sc_hd__a21oi_1
X_3604_ _3605_/B _3604_/B vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__and2b_1
X_3535_ _3536_/A _3536_/B _3536_/C vssd1 vssd1 vccd1 vccd1 _3535_/Y sky130_fd_sc_hd__a21oi_1
X_6323_ _6369_/CLK _6323_/D vssd1 vssd1 vccd1 vccd1 _6323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6254_ _6258_/C _6254_/B vssd1 vssd1 vccd1 vccd1 _6376_/D sky130_fd_sc_hd__nor2_1
X_3466_ _3465_/A _3465_/B _3465_/C vssd1 vssd1 vccd1 vccd1 _3471_/B sky130_fd_sc_hd__a21o_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5205_ _5469_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5489_/B sky130_fd_sc_hd__and2_2
X_6185_ _6344_/Q _6183_/X _6184_/X _6292_/D vssd1 vssd1 vccd1 vccd1 _6185_/X sky130_fd_sc_hd__o31a_1
X_3397_ _6304_/Q _6303_/Q _6296_/Q _6295_/Q _6294_/Q vssd1 vssd1 vccd1 vccd1 _3449_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5136_ _5136_/A _5136_/B _5215_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _5142_/A sky130_fd_sc_hd__or4bb_1
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5067_ _5273_/B vssd1 vssd1 vccd1 vccd1 _5388_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4018_/A _4018_/B vssd1 vssd1 vccd1 vccd1 _4018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3823__A1 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _5969_/A _5969_/B vssd1 vssd1 vccd1 vccd1 _5970_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5037__B _5059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3511__B1 _3536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_96 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3320_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3320_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3251_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3211__A _3214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5823_ _6382_/Q _5822_/X _5818_/Y _6383_/Q vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4230__A1 _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5754_ _6364_/Q _5713_/Y _5731_/Y _5732_/Y _5753_/X vssd1 vssd1 vccd1 vccd1 _5754_/X
+ sky130_fd_sc_hd__a2111o_1
X_4705_ _4705_/A _4705_/B vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__nor2_2
X_5685_ _5685_/A vssd1 vssd1 vccd1 vccd1 _5779_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4636_ _4701_/B _4636_/B vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4567_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5634_/A sky130_fd_sc_hd__buf_2
X_6306_ _6357_/CLK _6306_/D vssd1 vssd1 vccd1 vccd1 _6306_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5730__B2 _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4498_ _4484_/C _4488_/A _3924_/Y vssd1 vssd1 vccd1 vccd1 _4499_/D sky130_fd_sc_hd__a21o_1
X_3518_ _6295_/Q vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6237_ _6259_/A _6237_/B _6241_/C vssd1 vssd1 vccd1 vccd1 _6370_/D sky130_fd_sc_hd__nor3_1
X_3449_ _3449_/A _4814_/C vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__xnor2_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6343_/Q _6176_/B vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__and2_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5119_ _5119_/A _5550_/A vssd1 vssd1 vccd1 vccd1 _5120_/B sky130_fd_sc_hd__and2_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6099_ _6317_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6100_/A sky130_fd_sc_hd__and2_1
XFILLER_53_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6061__B _6061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5470_ _5470_/A _5476_/B vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__xnor2_1
X_4421_ _4421_/A _4421_/B vssd1 vssd1 vccd1 vccd1 _4423_/B sky130_fd_sc_hd__xnor2_1
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _4338_/A _4352_/B vssd1 vssd1 vccd1 vccd1 _4353_/B sky130_fd_sc_hd__and2b_1
X_4283_ _4284_/B _4283_/B vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3303_ _3306_/A vssd1 vssd1 vccd1 vccd1 _3303_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3206__A _3208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_577 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3234_ _3258_/A vssd1 vssd1 vccd1 vccd1 _3239_/A sky130_fd_sc_hd__buf_8
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6016_/A _5988_/X _6021_/X _6013_/X vssd1 vssd1 vccd1 vccd1 _6298_/D sky130_fd_sc_hd__o211a_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ _5386_/A vssd1 vssd1 vccd1 vccd1 _5314_/A sky130_fd_sc_hd__clkbuf_2
X_5806_ _5787_/Y _5790_/Y _5791_/Y _5802_/Y _5805_/Y vssd1 vssd1 vccd1 vccd1 _5806_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5737_ _5737_/A _5737_/B _5737_/C vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__and3_1
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5668_ _5583_/X _5584_/Y _5594_/X _5595_/X _5667_/X vssd1 vssd1 vccd1 vccd1 _5668_/X
+ sky130_fd_sc_hd__a2111o_1
X_4619_ _4619_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4619_/X sky130_fd_sc_hd__and2_1
X_5599_ _5737_/A _5652_/A vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__or2_1
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_634 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3953__B1 _5885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4970_ _5145_/B vssd1 vssd1 vccd1 vccd1 _4994_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3921_ _4479_/B _3968_/B vssd1 vssd1 vccd1 vccd1 _4492_/A sky130_fd_sc_hd__or2_1
XFILLER_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _5059_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__nand2_1
X_6571_ _6571_/A _3297_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_3783_ _3783_/A vssd1 vssd1 vccd1 vccd1 _3840_/A sky130_fd_sc_hd__clkbuf_2
X_5522_ _5522_/A _5521_/A vssd1 vssd1 vccd1 vccd1 _5523_/B sky130_fd_sc_hd__or2b_1
X_5453_ _5473_/A _5473_/B vssd1 vssd1 vccd1 vccd1 _5456_/B sky130_fd_sc_hd__and2_1
X_5384_ _5398_/A _5398_/B vssd1 vssd1 vccd1 vccd1 _5384_/X sky130_fd_sc_hd__and2_1
X_4404_ _4405_/A _4405_/B vssd1 vssd1 vccd1 vccd1 _4408_/B sky130_fd_sc_hd__xor2_1
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4335_ _4334_/A _4376_/B _4334_/C vssd1 vssd1 vccd1 vccd1 _4336_/B sky130_fd_sc_hd__a21oi_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_92 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4266_ _4266_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4274_/B sky130_fd_sc_hd__nand2_1
X_3217_ _3220_/A vssd1 vssd1 vccd1 vccd1 _3217_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4197_ _5450_/B _4412_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__nand2_1
X_6005_ _6000_/A _5988_/X _6004_/Y _5945_/X vssd1 vssd1 vccd1 vccd1 _6296_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5492__A1_N _4266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4120_ _5231_/A _4268_/B vssd1 vssd1 vccd1 vccd1 _4120_/X sky130_fd_sc_hd__and2_1
X_4051_ _4059_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4953_ _4953_/A _4953_/B vssd1 vssd1 vccd1 vccd1 _4954_/B sky130_fd_sc_hd__xor2_1
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3904_ _3950_/B vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _4731_/B _4864_/C _4714_/B _3631_/A vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__a22oi_1
X_3835_ _5274_/A vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6554_ _6554_/A _3267_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_3766_ _4634_/A _3502_/X _3734_/B _4698_/A vssd1 vssd1 vccd1 vccd1 _3768_/B sky130_fd_sc_hd__a22oi_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5505_ _5510_/A _5505_/B _5505_/C vssd1 vssd1 vccd1 vccd1 _5519_/A sky130_fd_sc_hd__and3_1
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3697_ _4814_/A _3697_/B _3697_/C _3503_/A vssd1 vssd1 vccd1 vccd1 _3739_/A sky130_fd_sc_hd__or4b_2
X_5436_ _6277_/Q _5291_/A _5439_/B _6278_/Q vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__a22o_1
XFILLER_105_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4985__A _5619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5367_ _6281_/Q _5394_/B _5439_/B vssd1 vssd1 vccd1 vccd1 _5367_/X sky130_fd_sc_hd__and3_1
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5298_ _5298_/A _5298_/B vssd1 vssd1 vccd1 vccd1 _5318_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4318_ _4346_/A _4346_/B _4316_/A vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__o21ai_1
X_4249_ _4250_/A _4250_/B vssd1 vssd1 vccd1 vccd1 _4251_/A sky130_fd_sc_hd__or2_1
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5312__C _5471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3304__A _3306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _3626_/A _3626_/B _3619_/Y vssd1 vssd1 vccd1 vccd1 _3624_/C sky130_fd_sc_hd__a21o_1
X_3551_ _4879_/B _3551_/B vssd1 vssd1 vccd1 vccd1 _3562_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3482_ _6287_/Q vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__inv_2
X_6270_ _6270_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _6270_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5221_ _5221_/A _5221_/B _5221_/C _5221_/D vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__nor4_2
X_5152_ _5113_/X _5149_/Y _5141_/X _5148_/X vssd1 vssd1 vccd1 vccd1 _5153_/C sky130_fd_sc_hd__a211o_1
XFILLER_69_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4103_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4477_/B sky130_fd_sc_hd__xnor2_2
XFILLER_96_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5413__B _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5083_ _5083_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _5552_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__3214__A _3214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4627__A1 _5702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ _4119_/A _4089_/A _3987_/B vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__or3b_1
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5985_ _6350_/Q _6359_/Q vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__and2b_1
X_4936_ _4953_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__and2b_1
XFILLER_52_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4867_ _4867_/A _4867_/B vssd1 vssd1 vccd1 vccd1 _4869_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3818_ _3818_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3840_/B sky130_fd_sc_hd__xnor2_2
X_4798_ _4798_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4800_/B sky130_fd_sc_hd__xor2_1
X_6537_ _6537_/A _3248_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3749_ _3749_/A _3749_/B vssd1 vssd1 vccd1 vccd1 _3782_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5419_ _5278_/A _5404_/B _5427_/A _5418_/X vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__a31o_1
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4519__B_N _4569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5993__B _6000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5034__B2 _5011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5770_ _5770_/A vssd1 vssd1 vccd1 vccd1 _6061_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4733_/C sky130_fd_sc_hd__nand2_1
X_6528__47 vssd1 vssd1 vccd1 vccd1 _6528__47/HI _6528_/A sky130_fd_sc_hd__conb_1
X_4652_ _4652_/A vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__buf_2
X_3603_ _3600_/Y _3632_/A _3602_/X _4882_/A vssd1 vssd1 vccd1 vccd1 _3604_/B sky130_fd_sc_hd__a2bb2o_1
X_4583_ _4583_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4583_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4312__B _6280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3534_ _3565_/A _3565_/B vssd1 vssd1 vccd1 vccd1 _3534_/Y sky130_fd_sc_hd__nand2_1
X_6322_ _6369_/CLK _6322_/D vssd1 vssd1 vccd1 vccd1 _6322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6253_ _6376_/Q vssd1 vssd1 vccd1 vccd1 _6258_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _3465_/A _3465_/B _3465_/C vssd1 vssd1 vccd1 vccd1 _3471_/A sky130_fd_sc_hd__nand3_1
X_5204_ _5203_/A _5203_/B _5203_/C vssd1 vssd1 vccd1 vccd1 _5469_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6184_ _6347_/Q _6346_/Q _6349_/Q _6348_/Q vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__or4_1
X_3396_ _6063_/A _6060_/A _5770_/A vssd1 vssd1 vccd1 vccd1 _3396_/Y sky130_fd_sc_hd__nor3_2
XFILLER_111_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5135_ _5134_/A _5134_/B _5134_/C vssd1 vssd1 vccd1 vccd1 _5136_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5066_ _5066_/A _5066_/B vssd1 vssd1 vccd1 vccd1 _5273_/B sky130_fd_sc_hd__xor2_4
X_4017_ _4017_/A _4017_/B vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__nor2_4
XANTENNA__3879__A _5646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _3379_/A _5949_/X _5967_/X vssd1 vssd1 vccd1 vccd1 _5969_/B sky130_fd_sc_hd__o21a_1
X_4919_ _5029_/A _5029_/B _4918_/Y vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5899_ _5899_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3250_/Y sky130_fd_sc_hd__inv_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4307__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5822_ _5698_/A _5820_/X _5821_/X _5706_/X vssd1 vssd1 vccd1 vccd1 _5822_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _6362_/Q _5734_/Y _5743_/X _5744_/X _5752_/X vssd1 vssd1 vccd1 vccd1 _5753_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4704_ _4704_/A _4743_/A _4704_/C vssd1 vssd1 vccd1 vccd1 _4705_/B sky130_fd_sc_hd__and3_1
X_5684_ _5703_/A _5759_/A _5675_/A vssd1 vssd1 vccd1 vccd1 _5684_/X sky130_fd_sc_hd__a21bo_1
X_4635_ _4634_/A _4931_/A _4638_/A vssd1 vssd1 vccd1 vccd1 _4636_/B sky130_fd_sc_hd__a21oi_1
X_4566_ _4566_/A _4566_/B vssd1 vssd1 vccd1 vccd1 _4569_/B sky130_fd_sc_hd__and2_1
XFILLER_116_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6305_ _6357_/CLK _6305_/D vssd1 vssd1 vccd1 vccd1 _6305_/Q sky130_fd_sc_hd__dfxtp_1
X_3517_ _3517_/A vssd1 vssd1 vccd1 vccd1 _5995_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4497_ _3937_/X _4492_/B _4490_/B _4491_/A vssd1 vssd1 vccd1 vccd1 _4499_/C sky130_fd_sc_hd__a211o_1
X_6236_ _6370_/Q _6369_/Q _6368_/Q vssd1 vssd1 vccd1 vccd1 _6241_/C sky130_fd_sc_hd__and3_1
X_3448_ _3405_/X _3406_/X _6297_/Q vssd1 vssd1 vccd1 vccd1 _4814_/C sky130_fd_sc_hd__a21oi_2
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6176_/B sky130_fd_sc_hd__clkbuf_1
X_3379_ _3379_/A _5957_/A vssd1 vssd1 vccd1 vccd1 _3380_/C sky130_fd_sc_hd__or2_1
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5118_ _5118_/A _5119_/A _5118_/C vssd1 vssd1 vccd1 vccd1 _5550_/A sky130_fd_sc_hd__nand3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6098_ _6098_/A vssd1 vssd1 vccd1 vccd1 _6107_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_84_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5049_ _5080_/A _5080_/B vssd1 vssd1 vccd1 vccd1 _5056_/C sky130_fd_sc_hd__and2b_1
XFILLER_27_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5064__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4857__B_N _4865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_654 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5511__B _5511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3312__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4420_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__inv_2
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4351_ _4354_/B _4354_/A vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__or2b_1
X_3302_ _3306_/A vssd1 vssd1 vccd1 vccd1 _3302_/Y sky130_fd_sc_hd__inv_2
X_4282_ _4194_/A _4370_/B _4280_/A _4311_/A vssd1 vssd1 vccd1 vccd1 _4283_/B sky130_fd_sc_hd__a31o_1
XFILLER_3_190 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3233_ input1/X vssd1 vssd1 vccd1 vccd1 _3258_/A sky130_fd_sc_hd__buf_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6019_/X _6026_/B _6023_/A vssd1 vssd1 vccd1 vccd1 _6021_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5702__A _5702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3222__A _3226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3997_ _4334_/A vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__clkbuf_2
X_5805_ _6372_/Q _5805_/B vssd1 vssd1 vccd1 vccd1 _5805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5736_ _5773_/A _5793_/A _5793_/B vssd1 vssd1 vccd1 vccd1 _5736_/X sky130_fd_sc_hd__or3_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _5601_/A _5593_/X _5599_/X _5601_/Y _5666_/X vssd1 vssd1 vccd1 vccd1 _5667_/X
+ sky130_fd_sc_hd__o221a_1
X_4618_ _4618_/A _4618_/B vssd1 vssd1 vccd1 vccd1 _4618_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4511__A_N _5702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5598_ _5598_/A _5598_/B vssd1 vssd1 vccd1 vccd1 _5652_/A sky130_fd_sc_hd__xnor2_2
X_6512__31 vssd1 vssd1 vccd1 vccd1 _6512__31/HI _6512_/A sky130_fd_sc_hd__conb_1
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4549_ _4548_/B _4548_/C _5605_/A vssd1 vssd1 vccd1 vccd1 _4550_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6219_ _6363_/Q _6221_/C _6218_/Y vssd1 vssd1 vccd1 vccd1 _6363_/D sky130_fd_sc_hd__o21a_1
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_646 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3953__A1 _3840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4138__A _4138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3977__A _4337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _4482_/A _3920_/B vssd1 vssd1 vccd1 vccd1 _3968_/B sky130_fd_sc_hd__or2_1
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3851_ _3851_/A _3851_/B vssd1 vssd1 vccd1 vccd1 _4088_/B sky130_fd_sc_hd__xnor2_4
XFILLER_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3782_ _3782_/A _3782_/B _3781_/X vssd1 vssd1 vccd1 vccd1 _3783_/A sky130_fd_sc_hd__or3b_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6570_ _6570_/A _3318_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
X_5521_ _5521_/A _5522_/A vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__or2b_1
XANTENNA__5697__A1 _3333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5452_ _5452_/A _5452_/B vssd1 vssd1 vccd1 vccd1 _5473_/B sky130_fd_sc_hd__xor2_1
X_5383_ _5383_/A _5383_/B vssd1 vssd1 vccd1 vccd1 _5398_/B sky130_fd_sc_hd__xor2_1
X_4403_ _4403_/A _4403_/B vssd1 vssd1 vccd1 vccd1 _4405_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5416__B _5444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3217__A _3220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4334_ _4334_/A _4334_/B _4334_/C vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__and3_1
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4265_ _4265_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__xnor2_1
X_6004_ _6057_/A _6004_/B vssd1 vssd1 vccd1 vccd1 _6004_/Y sky130_fd_sc_hd__nand2_1
X_4196_ _5394_/A vssd1 vssd1 vccd1 vccd1 _5450_/B sky130_fd_sc_hd__clkbuf_2
X_3216_ _3220_/A vssd1 vssd1 vccd1 vccd1 _3216_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4048__A _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5607__A _5675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5719_ _5719_/A _5719_/B vssd1 vssd1 vccd1 vccd1 _5719_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_21 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_484 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3797__A _4266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ _5236_/A vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput6 io_in[8] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4694_/B _4933_/B _4950_/Y _4951_/Y vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__a31o_1
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4883_ _4888_/A _4882_/C _4882_/A vssd1 vssd1 vccd1 vccd1 _4894_/B sky130_fd_sc_hd__o21ai_1
X_3834_ _5381_/A vssd1 vssd1 vccd1 vccd1 _5274_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3765_ _3805_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__xnor2_1
X_6553_ _6553_/A _3263_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_3696_ _3696_/A _3696_/B vssd1 vssd1 vccd1 vccd1 _3697_/B sky130_fd_sc_hd__nand2_1
X_5504_ _5504_/A _5504_/B vssd1 vssd1 vccd1 vccd1 _5520_/B sky130_fd_sc_hd__or2_1
X_5435_ _5435_/A _5435_/B vssd1 vssd1 vccd1 vccd1 _5533_/A sky130_fd_sc_hd__xnor2_2
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _5324_/A _5439_/B _4280_/B vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__a21bo_1
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5297_ _5297_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5298_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5162__A _5382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4317_ _4317_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4346_/B sky130_fd_sc_hd__xnor2_1
X_4248_ _4276_/A _4275_/B _4275_/A vssd1 vssd1 vccd1 vccd1 _4250_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4179_ _4141_/C _4142_/X _4175_/X _4181_/A vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__a211oi_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4225__B _4396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3320__A _3321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3550_ _6284_/Q vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5214_/A _5214_/B _5213_/X vssd1 vssd1 vccd1 vccd1 _5221_/D sky130_fd_sc_hd__o21ba_1
X_6588__104 vssd1 vssd1 vccd1 vccd1 _6588__104/HI _6588_/A sky130_fd_sc_hd__conb_1
X_3481_ _6291_/Q vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__inv_2
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5151_ _5151_/A _5151_/B vssd1 vssd1 vccd1 vccd1 _5153_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4102_ _4100_/A _4100_/B _4101_/X vssd1 vssd1 vccd1 vccd1 _4477_/A sky130_fd_sc_hd__a21o_2
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5082_ _5082_/A _5554_/C vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__5413__C _5469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4033_ _3782_/A _3720_/B _5885_/A vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__a21o_1
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5710__A _5710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3230__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5984_ _6359_/Q _6350_/Q vssd1 vssd1 vccd1 vccd1 _5984_/X sky130_fd_sc_hd__and2b_1
X_4935_ _4933_/A _4933_/B _4933_/D _4934_/X vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__a22o_1
X_4866_ _4898_/B _4866_/B vssd1 vssd1 vccd1 vccd1 _4867_/B sky130_fd_sc_hd__nor2_1
X_3817_ _3781_/A _3781_/B _3778_/A vssd1 vssd1 vccd1 vccd1 _3818_/B sky130_fd_sc_hd__a21o_1
X_4797_ _4797_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4798_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6554__70 vssd1 vssd1 vccd1 vccd1 _6554__70/HI _6554_/A sky130_fd_sc_hd__conb_1
XANTENNA__4061__A _4138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ _3717_/A _3717_/B _3717_/C _3715_/A vssd1 vssd1 vccd1 vccd1 _3749_/B sky130_fd_sc_hd__a31o_1
X_6536_ _6536_/A _3247_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_3679_ _5324_/A vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5418_ _5418_/A _5418_/B vssd1 vssd1 vccd1 vccd1 _5418_/X sky130_fd_sc_hd__and2_1
XFILLER_99_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5349_ _5349_/A _5444_/B _5444_/C vssd1 vssd1 vccd1 vccd1 _5362_/B sky130_fd_sc_hd__and3_1
XFILLER_102_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5620__A _5627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5067__A _5273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3315__A _3318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4146__A _5246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4733_/B _4720_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__and2_1
XFILLER_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5990__B1 _5952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4651_ _4651_/A vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__inv_2
X_3602_ _4864_/B _3600_/B _3601_/B _4842_/B vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__a22o_1
X_4582_ _4583_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4586_/B sky130_fd_sc_hd__xor2_1
XFILLER_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3533_ _3540_/A _3540_/B vssd1 vssd1 vccd1 vccd1 _3565_/B sky130_fd_sc_hd__xor2_1
X_6321_ _6369_/CLK _6321_/D vssd1 vssd1 vccd1 vccd1 _6321_/Q sky130_fd_sc_hd__dfxtp_1
X_6252_ _6375_/Q _6249_/B _6251_/Y vssd1 vssd1 vccd1 vccd1 _6375_/D sky130_fd_sc_hd__o21a_1
X_3464_ _3464_/A _3464_/B vssd1 vssd1 vccd1 vccd1 _3465_/C sky130_fd_sc_hd__xor2_1
XFILLER_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _5203_/A _5203_/B _5203_/C vssd1 vssd1 vccd1 vccd1 _5469_/B sky130_fd_sc_hd__nand3_2
X_6183_ _6343_/Q _6342_/Q _6345_/Q vssd1 vssd1 vccd1 vccd1 _6183_/X sky130_fd_sc_hd__or3_1
X_5134_ _5134_/A _5134_/B _5134_/C vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__and3_1
XANTENNA__3225__A _3226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3395_ _5814_/C vssd1 vssd1 vccd1 vccd1 _5770_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5065_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _5074_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4016_ _4016_/A _4016_/B _4016_/C vssd1 vssd1 vccd1 vccd1 _4017_/B sky130_fd_sc_hd__and3_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ _3380_/C _5966_/B _5959_/X vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _4918_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _4918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5898_ _5898_/A vssd1 vssd1 vccd1 vccd1 _6278_/D sky130_fd_sc_hd__clkbuf_1
X_4849_ _4844_/B _4866_/B _4844_/A vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__a21bo_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6519_ _6519_/A _3226_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_106_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5615__A _5672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3789__B _3947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5821_ _5690_/B _5702_/Y _5703_/Y _5773_/B vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__o22a_1
X_5752_ _6361_/Q _5739_/X _5741_/Y _5751_/Y _6360_/Q vssd1 vssd1 vccd1 vccd1 _5752_/X
+ sky130_fd_sc_hd__a311o_1
X_4703_ _4704_/A _4743_/A _4704_/C vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5683_ _5683_/A _5683_/B _5711_/B vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__and3_1
X_4634_ _4634_/A _4931_/A _4638_/A vssd1 vssd1 vccd1 vccd1 _4701_/B sky130_fd_sc_hd__and3_1
X_4565_ _4565_/A _4565_/B vssd1 vssd1 vccd1 vccd1 _4566_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4034__C_N _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6304_ _6335_/CLK _6304_/D vssd1 vssd1 vccd1 vccd1 _6304_/Q sky130_fd_sc_hd__dfxtp_1
X_3516_ _3516_/A _3645_/C vssd1 vssd1 vccd1 vccd1 _3516_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4496_ _4496_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__or2_1
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235_ _5801_/A _6232_/A _6370_/Q vssd1 vssd1 vccd1 vccd1 _6237_/B sky130_fd_sc_hd__a21oi_1
X_3447_ _6290_/Q _3559_/B _3446_/C _3446_/D vssd1 vssd1 vccd1 vccd1 _3452_/B sky130_fd_sc_hd__a22o_1
XANTENNA__6291__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3378_ _4634_/A vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__buf_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5117_ _5114_/X _5115_/Y _5106_/Y _5113_/X vssd1 vssd1 vccd1 vccd1 _5118_/C sky130_fd_sc_hd__o211ai_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6097_ _6097_/A vssd1 vssd1 vccd1 vccd1 _6317_/D sky130_fd_sc_hd__clkbuf_1
X_5048_ _5056_/B _5048_/B vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_416 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4514__A _4555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_64 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__xor2_1
X_3301_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3306_/A sky130_fd_sc_hd__clkbuf_8
X_4281_ _5394_/A _4389_/A _4281_/C vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__and3_1
X_3232_ _3232_/A vssd1 vssd1 vccd1 vccd1 _3232_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _6020_/A _6020_/B vssd1 vssd1 vccd1 vccd1 _6026_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5804_ _5890_/A _5778_/X _5803_/X _3384_/X vssd1 vssd1 vccd1 vccd1 _5805_/B sky130_fd_sc_hd__a22oi_1
XANTENNA__4334__A _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3996_ _5485_/A vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4053__B _4088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5735_ _5735_/A _5735_/B _5747_/A vssd1 vssd1 vccd1 vccd1 _5793_/B sky130_fd_sc_hd__and3_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3962__A2 _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5666_ _5599_/X _5601_/Y _5612_/X _5665_/X vssd1 vssd1 vccd1 vccd1 _5666_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4617_ _4511_/X _4617_/B vssd1 vssd1 vccd1 vccd1 _4617_/X sky130_fd_sc_hd__and2b_1
X_5597_ _5597_/A _5597_/B vssd1 vssd1 vccd1 vccd1 _5737_/A sky130_fd_sc_hd__xnor2_4
X_4548_ _4548_/A _4548_/B _4548_/C vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__and3_1
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4479_ _4479_/A _4479_/B _4479_/C vssd1 vssd1 vccd1 vccd1 _4521_/B sky130_fd_sc_hd__and3_1
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6218_ _6218_/A _6218_/B vssd1 vssd1 vccd1 vccd1 _6218_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6149_ _6336_/Q _6165_/B vssd1 vssd1 vccd1 vccd1 _6150_/A sky130_fd_sc_hd__and2_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4228__B _4337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5059__B _5059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3953__A2 _3785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4898__B _4898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4138__B _4138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3977__B _4337_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _5098_/A vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6186__A3 _5861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3781_ _3781_/A _3781_/B vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__xor2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5520_ _5520_/A _5520_/B vssd1 vssd1 vccd1 vccd1 _5522_/A sky130_fd_sc_hd__xor2_1
X_5451_ _5451_/A _5451_/B vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__or2_1
X_5382_ _5382_/A _5382_/B _5382_/C vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__and3_1
X_4402_ _4421_/A _4421_/B vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5416__C _5444_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4333_ _5382_/A _4340_/B _4330_/X _4332_/Y vssd1 vssd1 vccd1 vccd1 _4334_/C sky130_fd_sc_hd__a31o_1
XFILLER_101_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4264_ _5381_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__and2_1
XFILLER_113_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3215_ _3227_/A vssd1 vssd1 vccd1 vccd1 _3220_/A sky130_fd_sc_hd__buf_8
X_6003_ _6003_/A _6003_/B vssd1 vssd1 vccd1 vccd1 _6004_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3233__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4195_ _6279_/Q vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3887__B _4166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _5166_/A _4323_/B vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__nand2_1
X_5718_ _5574_/Y _5678_/X _5680_/Y _5681_/Y vssd1 vssd1 vccd1 vccd1 _5719_/B sky130_fd_sc_hd__o211a_1
XFILLER_6_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4511__B _4555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5649_ _5652_/A _5652_/B vssd1 vssd1 vccd1 vccd1 _5651_/B sky130_fd_sc_hd__or2_1
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5623__A _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3318__A _3318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6352__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput7 io_in[9] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_36_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4951_ _3380_/A _4933_/B _4950_/Y _4694_/B vssd1 vssd1 vccd1 vccd1 _4951_/Y sky130_fd_sc_hd__a22oi_1
X_3902_ _3902_/A _3902_/B vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__nor2_1
X_4882_ _4882_/A _4888_/A _4882_/C vssd1 vssd1 vccd1 vccd1 _4894_/A sky130_fd_sc_hd__or3_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3833_ _5440_/A vssd1 vssd1 vccd1 vccd1 _5381_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3764_ _3764_/A _3764_/B vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__xnor2_1
X_6552_ _6552_/A _3261_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_5503_ _4266_/A _5510_/B _5484_/B vssd1 vssd1 vccd1 vccd1 _5504_/B sky130_fd_sc_hd__a21oi_1
X_3695_ _3647_/A _3647_/C _3647_/B vssd1 vssd1 vccd1 vccd1 _3702_/A sky130_fd_sc_hd__o21bai_1
X_5434_ _5535_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5598_/A sky130_fd_sc_hd__xor2_2
XANTENNA__3228__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5365_ _5505_/B vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__clkbuf_2
X_5296_ _5297_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5298_/A sky130_fd_sc_hd__or2_1
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4316_ _4316_/A _4316_/B vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4059__A _4059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4247_ _5328_/A _4361_/B _4280_/A vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__and3_1
X_4178_ _4180_/A _4180_/B _4180_/C vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__o21a_1
XFILLER_74_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4333__A2 _4340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3601__A _3601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3480_ _3645_/C vssd1 vssd1 vccd1 vccd1 _3600_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5150_ _5141_/X _5148_/X _5113_/X _5149_/Y vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__o211ai_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4101_ _4105_/A _4105_/B vssd1 vssd1 vccd1 vccd1 _4101_/X sky130_fd_sc_hd__and2_1
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5081_ _5083_/B _5083_/A vssd1 vssd1 vccd1 vccd1 _5554_/C sky130_fd_sc_hd__and2b_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _5231_/A vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__inv_2
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5983_ _6292_/Q _6313_/Q vssd1 vssd1 vccd1 vccd1 _5983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4934_ _5966_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__or2_1
X_4865_ _4865_/A _4885_/A vssd1 vssd1 vccd1 vccd1 _4867_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3816_ _3816_/A _3816_/B vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__and2_1
X_4796_ _4796_/A _4864_/B _4820_/B _4796_/D vssd1 vssd1 vccd1 vccd1 _4797_/B sky130_fd_sc_hd__and4_1
X_3747_ _3747_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__nor2_1
X_6535_ _6535_/A _3245_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5061__D_N _5038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3678_ _6280_/Q vssd1 vssd1 vccd1 vccd1 _5324_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5417_ _5418_/A _5418_/B vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__xor2_2
X_5348_ _4331_/A _5471_/B _5471_/C _5489_/B _5381_/A vssd1 vssd1 vccd1 vccd1 _5348_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_101_132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5279_ _5300_/A _5300_/B vssd1 vssd1 vccd1 vccd1 _5279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5901__A _5901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5503__A1 _4266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4146__B _4396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _4680_/A _4680_/B _4648_/X vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3601_ _3601_/A _3601_/B vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__nand2_1
X_4581_ _4581_/A _4581_/B vssd1 vssd1 vccd1 vccd1 _4583_/B sky130_fd_sc_hd__xor2_1
X_6320_ _6369_/CLK _6320_/D vssd1 vssd1 vccd1 vccd1 _6320_/Q sky130_fd_sc_hd__dfxtp_1
X_3532_ _3532_/A _3532_/B vssd1 vssd1 vccd1 vccd1 _3540_/B sky130_fd_sc_hd__xor2_1
X_6251_ _6375_/Q _6249_/B _6218_/A vssd1 vssd1 vccd1 vccd1 _6251_/Y sky130_fd_sc_hd__a21oi_1
X_3463_ _3463_/A _3463_/B vssd1 vssd1 vccd1 vccd1 _3464_/B sky130_fd_sc_hd__or2_1
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5202_ _5202_/A _5202_/B vssd1 vssd1 vccd1 vccd1 _5211_/A sky130_fd_sc_hd__xnor2_1
X_6182_ _6342_/Q _6345_/Q _6182_/C vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__and3_1
X_5133_ _5133_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5134_/C sky130_fd_sc_hd__and2_1
X_3394_ _6302_/Q vssd1 vssd1 vccd1 vccd1 _5814_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5064_ _5064_/A _5180_/D vssd1 vssd1 vccd1 vccd1 _5065_/A sky130_fd_sc_hd__nand2_1
X_4015_ _4016_/A _4016_/B _4016_/C vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__3241__A _3245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5966_ _5966_/A _5966_/B vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__xnor2_1
X_4917_ _5066_/A _5066_/B _4916_/X vssd1 vssd1 vccd1 vccd1 _5029_/B sky130_fd_sc_hd__a21o_2
X_5897_ _6140_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5898_/A sky130_fd_sc_hd__and2_1
X_4848_ _4852_/C _4852_/B _4869_/A vssd1 vssd1 vccd1 vccd1 _4854_/A sky130_fd_sc_hd__a21bo_1
X_6519__38 vssd1 vssd1 vccd1 vccd1 _6519__38/HI _6519_/A sky130_fd_sc_hd__conb_1
XFILLER_20_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4779_ _4778_/B _4779_/B vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__and2b_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4800__A _4818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6518_ _6518_/A _3225_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_506 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5350__B _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6533__52 vssd1 vssd1 vccd1 vccd1 _6533__52/HI _6533_/A sky130_fd_sc_hd__conb_1
XFILLER_98_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5820_ _5820_/A vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5751_ _5867_/A _5741_/B _5750_/X _3383_/A vssd1 vssd1 vccd1 vccd1 _5751_/Y sky130_fd_sc_hd__a22oi_1
X_4702_ _4941_/A _4702_/B vssd1 vssd1 vccd1 vccd1 _4704_/C sky130_fd_sc_hd__nor2_1
X_5682_ _5574_/Y _5678_/X _5719_/A _5680_/Y _5681_/Y vssd1 vssd1 vccd1 vccd1 _5711_/B
+ sky130_fd_sc_hd__o2111a_1
X_4633_ _4731_/A _4694_/A _4714_/B _4846_/B vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__and4_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ _5627_/A _4564_/B vssd1 vssd1 vccd1 vccd1 _4564_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6303_ _6335_/CLK _6303_/D vssd1 vssd1 vccd1 vccd1 _6303_/Q sky130_fd_sc_hd__dfxtp_1
X_3515_ _3515_/A _3515_/B vssd1 vssd1 vccd1 vccd1 _3527_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3236__A _3239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4495_ _4495_/A _4495_/B vssd1 vssd1 vccd1 vccd1 _5710_/A sky130_fd_sc_hd__xor2_4
X_6234_ _5801_/A _6232_/A _6233_/Y vssd1 vssd1 vccd1 vccd1 _6369_/D sky130_fd_sc_hd__o21a_1
X_3446_ _4651_/A _3601_/B _3446_/C _3446_/D vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__nand4_1
X_3377_ _3377_/A vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__clkbuf_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6342_/Q _6165_/B vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__and2_1
X_5116_ _5106_/Y _5113_/X _5114_/X _5115_/Y vssd1 vssd1 vccd1 vccd1 _5119_/A sky130_fd_sc_hd__a211o_1
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6096_ _6316_/Q _6096_/B vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__and2_1
X_5047_ _5047_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5048_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5954__A1 _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5949_ _5966_/B vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4514__B _5702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6309__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5255__B _5358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3300_/Y sky130_fd_sc_hd__inv_2
X_4280_ _4280_/A _4280_/B vssd1 vssd1 vccd1 vccd1 _4281_/C sky130_fd_sc_hd__xnor2_1
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3231_ _3232_/A vssd1 vssd1 vccd1 vccd1 _3231_/Y sky130_fd_sc_hd__inv_2
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5803_ _5769_/X _5711_/Y _5771_/Y _5710_/X vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__a22o_1
X_3995_ _6275_/Q vssd1 vssd1 vccd1 vccd1 _5485_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _3384_/A _5728_/X _5700_/X _5733_/X vssd1 vssd1 vccd1 vccd1 _5734_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__3411__A2 _4814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5665_ _5612_/A _5610_/X _5618_/Y _5663_/X _5664_/Y vssd1 vssd1 vccd1 vccd1 _5665_/X
+ sky130_fd_sc_hd__a221o_1
X_4616_ _4542_/X _4612_/X _4614_/X _4615_/Y vssd1 vssd1 vccd1 vccd1 _4616_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5165__B _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5596_ _5550_/X _5596_/B vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__and2b_1
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ _4546_/A _4546_/B _4546_/C vssd1 vssd1 vccd1 vccd1 _4548_/C sky130_fd_sc_hd__a21o_1
X_4478_ _4506_/A _4506_/B _4531_/A _4477_/X vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__a211o_1
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3429_ _4846_/A _3503_/A _3503_/B vssd1 vssd1 vccd1 vccd1 _3473_/A sky130_fd_sc_hd__and3_1
X_6217_ _6363_/Q _6221_/C vssd1 vssd1 vccd1 vccd1 _6218_/B sky130_fd_sc_hd__and2_1
XFILLER_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6148_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6165_/B sky130_fd_sc_hd__clkbuf_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4228__C _4337_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _6079_/A vssd1 vssd1 vccd1 vccd1 _6311_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4525__A _5710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6503__22 vssd1 vssd1 vccd1 vccd1 _6503__22/HI _6503_/A sky130_fd_sc_hd__conb_1
XFILLER_107_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6187__A _6187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5091__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3780_ _3717_/A _3717_/B _3717_/C _3749_/A _3779_/X vssd1 vssd1 vccd1 vccd1 _3781_/B
+ sky130_fd_sc_hd__a41o_1
X_5450_ _5936_/A _5450_/B _5450_/C vssd1 vssd1 vccd1 vccd1 _5473_/A sky130_fd_sc_hd__and3_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5146__A2 _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4401_ _4401_/A vssd1 vssd1 vccd1 vccd1 _4421_/B sky130_fd_sc_hd__inv_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5381_ _5381_/A _5486_/B vssd1 vssd1 vccd1 vccd1 _5383_/B sky130_fd_sc_hd__and2_1
XFILLER_5_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _4332_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ _4331_/A _4365_/B _4365_/C vssd1 vssd1 vccd1 vccd1 _4265_/A sky130_fd_sc_hd__and3_1
XFILLER_59_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3214_ _3214_/A vssd1 vssd1 vccd1 vccd1 _3214_/Y sky130_fd_sc_hd__inv_2
X_6002_ _5993_/A _6016_/B _5994_/X vssd1 vssd1 vccd1 vccd1 _6003_/B sky130_fd_sc_hd__a21oi_1
X_4194_ _4194_/A _4389_/A vssd1 vssd1 vccd1 vccd1 _4198_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3978_ _4076_/B vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5717_ _5717_/A _5717_/B vssd1 vssd1 vccd1 vccd1 _5717_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_109_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5648_ _5648_/A _5648_/B vssd1 vssd1 vccd1 vccd1 _5652_/B sky130_fd_sc_hd__nand2_1
X_5579_ _5579_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _5580_/B sky130_fd_sc_hd__nand2_2
XFILLER_2_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3424__A _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5073__B2 _5038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6575__91 vssd1 vssd1 vccd1 vccd1 _6575__91/HI _6575_/A sky130_fd_sc_hd__conb_1
XFILLER_107_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput8 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4950_ _5966_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3901_ _3901_/A _3894_/B vssd1 vssd1 vccd1 vccd1 _3916_/B sky130_fd_sc_hd__or2b_1
X_4881_ _4881_/A _4881_/B _4897_/A vssd1 vssd1 vccd1 vccd1 _4882_/C sky130_fd_sc_hd__and3_1
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _6278_/Q vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6551_ _6551_/A _3259_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3763_ _3763_/A _3807_/B vssd1 vssd1 vccd1 vccd1 _3764_/B sky130_fd_sc_hd__nand2_2
X_5502_ _5471_/A _5485_/B _5365_/X _5416_/A vssd1 vssd1 vccd1 vccd1 _5519_/B sky130_fd_sc_hd__a22oi_1
X_3694_ _3661_/A _3697_/C _3691_/X _3743_/A vssd1 vssd1 vccd1 vccd1 _3704_/A sky130_fd_sc_hd__a22o_1
X_5433_ _5435_/A _5435_/B _5432_/X vssd1 vssd1 vccd1 vccd1 _5535_/B sky130_fd_sc_hd__a21bo_1
X_5364_ _5370_/A _5370_/B vssd1 vssd1 vccd1 vccd1 _5369_/A sky130_fd_sc_hd__or2_1
XANTENNA__5724__A _5724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4315_ _4315_/A _4344_/A vssd1 vssd1 vccd1 vccd1 _4316_/B sky130_fd_sc_hd__or2_1
X_5295_ _5323_/A _5322_/B _5322_/A vssd1 vssd1 vccd1 vccd1 _5297_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3244__A _3245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6494__13 vssd1 vssd1 vccd1 vccd1 _6494__13/HI _6494_/A sky130_fd_sc_hd__conb_1
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4246_ _6280_/Q _4388_/B vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__and2_1
X_4177_ _4177_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4180_/C sky130_fd_sc_hd__xnor2_1
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5634__A _5634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5781__A1_N _5698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5263__B _5267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4100_ _4100_/A _4100_/B vssd1 vssd1 vccd1 vccd1 _4105_/B sky130_fd_sc_hd__xor2_1
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _5080_/A _5080_/B vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__xnor2_1
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4031_ _4031_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3999__A _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_275 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5982_ _6292_/Q _6313_/Q vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__and2_1
X_4933_ _4933_/A _4933_/B _4950_/B _4933_/D vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__and4_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4864_ _4879_/A _4864_/B _4864_/C _4864_/D vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__and4_1
XFILLER_20_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3815_ _3815_/A _3815_/B vssd1 vssd1 vccd1 vccd1 _3816_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5438__B _5486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _4791_/A _4791_/B _4788_/X vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__a21bo_1
X_3746_ _3746_/A _3746_/B vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__and2_1
X_6534_ _6534_/A _3244_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XANTENNA__3239__A _3239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3677_ _3940_/B vssd1 vssd1 vccd1 vccd1 _4168_/B sky130_fd_sc_hd__clkbuf_2
X_5416_ _5416_/A _5444_/B _5444_/C vssd1 vssd1 vccd1 vccd1 _5418_/B sky130_fd_sc_hd__and3_1
XFILLER_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5347_ _5347_/A _5347_/B vssd1 vssd1 vccd1 vccd1 _5539_/B sky130_fd_sc_hd__xnor2_4
X_5278_ _5278_/A _5278_/B vssd1 vssd1 vccd1 vccd1 _5300_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4229_ _4238_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__and2_1
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6545__61 vssd1 vssd1 vccd1 vccd1 _6545__61/HI _6545_/A sky130_fd_sc_hd__conb_1
XFILLER_7_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594__110 vssd1 vssd1 vccd1 vccd1 _6594__110/HI _6594_/A sky130_fd_sc_hd__conb_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4580_ _5183_/A _4580_/B _4587_/B vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__and3_1
X_3600_ _4785_/A _3600_/B vssd1 vssd1 vccd1 vccd1 _3600_/Y sky130_fd_sc_hd__nand2_1
X_3531_ _4879_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3532_/B sky130_fd_sc_hd__nand2_1
X_6250_ _6374_/Q _6246_/B _6249_/Y vssd1 vssd1 vccd1 vccd1 _6374_/D sky130_fd_sc_hd__o21a_1
X_3462_ _3520_/B _3479_/A _3522_/B _3494_/A vssd1 vssd1 vccd1 vccd1 _3463_/B sky130_fd_sc_hd__a22oi_1
X_5201_ _5243_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _5202_/A sky130_fd_sc_hd__nand2_1
X_6181_ _6347_/Q _6346_/Q _6349_/Q _6348_/Q vssd1 vssd1 vccd1 vccd1 _6182_/C sky130_fd_sc_hd__and4_1
X_3393_ _5701_/B vssd1 vssd1 vccd1 vccd1 _6060_/A sky130_fd_sc_hd__clkbuf_2
X_5132_ _5085_/A _5158_/B _5159_/B _5130_/X vssd1 vssd1 vccd1 vccd1 _5138_/B sky130_fd_sc_hd__a31o_1
XFILLER_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _5046_/B _5043_/B _5043_/C vssd1 vssd1 vccd1 vccd1 _5078_/B sky130_fd_sc_hd__a21oi_1
X_4014_ _4014_/A _4014_/B vssd1 vssd1 vccd1 vccd1 _4016_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__4337__B _4337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5965_ _3379_/A _5963_/X _5964_/Y vssd1 vssd1 vccd1 vccd1 _6289_/D sky130_fd_sc_hd__o21a_1
X_4916_ _4837_/B _4916_/B vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__and2b_1
XFILLER_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5896_ _5890_/A _5895_/Y _5896_/S vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__mux2_1
X_4847_ _4868_/B _4868_/C _4868_/A vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4778_ _4779_/B _4778_/B vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__xnor2_4
XFILLER_20_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6517_ _6517_/A _3224_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
X_3729_ _3729_/A _3729_/B vssd1 vssd1 vccd1 vccd1 _3746_/A sky130_fd_sc_hd__nand2_1
X_6379_ _6383_/CLK _6379_/D vssd1 vssd1 vccd1 vccd1 _6379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5350__C _5469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_448 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5541__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _3396_/Y _5747_/X _5749_/Y _5687_/X vssd1 vssd1 vccd1 vccd1 _5750_/X sky130_fd_sc_hd__a22o_1
X_4701_ _4701_/A _4701_/B _4701_/C vssd1 vssd1 vccd1 vccd1 _4702_/B sky130_fd_sc_hd__nor3_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _5737_/A vssd1 vssd1 vccd1 vccd1 _5681_/Y sky130_fd_sc_hd__inv_2
X_4632_ _4769_/B vssd1 vssd1 vccd1 vccd1 _4846_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4563_ _5619_/A _4563_/B vssd1 vssd1 vccd1 vccd1 _4563_/Y sky130_fd_sc_hd__xnor2_1
X_4494_ _4521_/A _4494_/B vssd1 vssd1 vccd1 vccd1 _4495_/B sky130_fd_sc_hd__nor2_2
X_6302_ _6359_/CLK _6302_/D vssd1 vssd1 vccd1 vccd1 _6302_/Q sky130_fd_sc_hd__dfxtp_1
X_3514_ _3514_/A _3514_/B vssd1 vssd1 vccd1 vccd1 _3515_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6233_ _5801_/A _6232_/A _6218_/A vssd1 vssd1 vccd1 vccd1 _6233_/Y sky130_fd_sc_hd__a21oi_1
X_3445_ _3516_/A _3549_/B _3549_/C _4877_/D _6291_/Q vssd1 vssd1 vccd1 vccd1 _3446_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3376_ _4645_/A vssd1 vssd1 vccd1 vccd1 _3377_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6164_/A vssd1 vssd1 vccd1 vccd1 _6342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5115_ _5114_/A _5114_/C _5114_/B vssd1 vssd1 vccd1 vccd1 _5115_/Y sky130_fd_sc_hd__a21oi_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6095_/A vssd1 vssd1 vccd1 vccd1 _6316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5046_ _5040_/A _5046_/B vssd1 vssd1 vccd1 vccd1 _5080_/A sky130_fd_sc_hd__and2b_1
XFILLER_27_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5948_ _5940_/A _3381_/B _5937_/A _5966_/B vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__a31o_1
XFILLER_43_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _5879_/A _5879_/B vssd1 vssd1 vccd1 vccd1 _5880_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3230_ _3232_/A vssd1 vssd1 vccd1 vccd1 _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5271__B _5444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_484 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5881__A1 _5733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_543 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5802_ _6371_/Q _5787_/B _5795_/X _5800_/X _5801_/X vssd1 vssd1 vccd1 vccd1 _5802_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3994_ _3994_/A _3994_/B vssd1 vssd1 vccd1 vccd1 _4005_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5733_ _5875_/A vssd1 vssd1 vccd1 vccd1 _5733_/X sky130_fd_sc_hd__clkbuf_2
X_5664_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5664_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4615_ _4615_/A _4615_/B vssd1 vssd1 vccd1 vccd1 _4615_/Y sky130_fd_sc_hd__nor2_1
X_5595_ _5669_/A _5669_/B vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__and2_1
XANTENNA__5165__C _5471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ _4546_/A _4546_/B _4546_/C vssd1 vssd1 vccd1 vccd1 _4548_/B sky130_fd_sc_hd__nand3_1
XANTENNA__3247__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4477_ _4477_/A _4477_/B vssd1 vssd1 vccd1 vccd1 _4477_/X sky130_fd_sc_hd__and2_1
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3428_ _6040_/A _3653_/B _4707_/B vssd1 vssd1 vccd1 vccd1 _3503_/B sky130_fd_sc_hd__or3_2
X_6216_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6218_/A sky130_fd_sc_hd__clkbuf_2
X_3359_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6147_ _6147_/A vssd1 vssd1 vccd1 vccd1 _6336_/D sky130_fd_sc_hd__clkbuf_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6078_ _6310_/Q _6096_/B vssd1 vssd1 vccd1 vccd1 _6079_/A sky130_fd_sc_hd__and2_1
X_5029_ _5029_/A _5029_/B vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__xor2_4
XANTENNA__4525__B _4569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5637__A _5637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6187__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _4400_/A _4400_/B vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5380_ _5380_/A _5380_/B vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4331_ _4331_/A _4361_/B vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4331_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__nand2_1
X_3213_ _3214_/A vssd1 vssd1 vccd1 vccd1 _3213_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6001_ _6001_/A _6001_/B vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _4361_/B vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4626__A _4626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3530__A _6285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3977_ _4337_/B _4337_/C vssd1 vssd1 vccd1 vccd1 _4076_/B sky130_fd_sc_hd__and2_1
X_5716_ _5735_/B _5747_/A _5724_/A _5735_/A vssd1 vssd1 vccd1 vccd1 _5717_/B sky130_fd_sc_hd__a211o_1
XFILLER_109_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _4138_/A _5510_/B _4587_/B vssd1 vssd1 vccd1 vccd1 _5648_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5578_ _5578_/A _5578_/B _5578_/C vssd1 vssd1 vccd1 vccd1 _5579_/B sky130_fd_sc_hd__or3_1
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4529_ _4624_/A _4577_/A vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6022__A1 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4033__B1 _5885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4584__A1 _5646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5367__A _6281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5814__B _6060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3900_ _3900_/A _3895_/A vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__or2b_1
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4880_ _4881_/A _4881_/B _4897_/A vssd1 vssd1 vccd1 vccd1 _4888_/A sky130_fd_sc_hd__a21oi_1
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3831_ _3877_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3762_ _4731_/A _3762_/B vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__nand2_1
X_6550_ _6550_/A _3256_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_9_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5501_ _5501_/A _5501_/B vssd1 vssd1 vccd1 vccd1 _5508_/A sky130_fd_sc_hd__xnor2_1
X_3693_ _3693_/A _3734_/C vssd1 vssd1 vccd1 vccd1 _3743_/A sky130_fd_sc_hd__nand2_1
X_5432_ _5432_/A _5431_/A vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__or2b_1
XFILLER_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5363_ _5450_/B _5485_/B _5330_/C vssd1 vssd1 vccd1 vccd1 _5370_/B sky130_fd_sc_hd__a21oi_1
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4314_ _4315_/A _4344_/A vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__nand2_1
XFILLER_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5294_ _5294_/A _5294_/B _5505_/B vssd1 vssd1 vccd1 vccd1 _5322_/A sky130_fd_sc_hd__and3_1
XANTENNA__5827__B2 _5733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4245_ _5324_/A _4389_/A _4409_/B _5328_/A vssd1 vssd1 vccd1 vccd1 _4275_/B sky130_fd_sc_hd__a22oi_1
X_4176_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4180_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3260__A _3263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5818__A1 _3333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4266__A _4266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3345__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _3981_/B _4075_/A _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4031_/B sky130_fd_sc_hd__o22ai_2
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5981_ _5981_/A vssd1 vssd1 vccd1 vccd1 _6293_/D sky130_fd_sc_hd__clkbuf_1
X_4932_ _4692_/A _4694_/B _4656_/A vssd1 vssd1 vccd1 vccd1 _4933_/D sky130_fd_sc_hd__a21bo_1
XFILLER_52_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4863_ _4854_/A _4853_/C _4853_/B vssd1 vssd1 vccd1 vccd1 _4870_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3814_ _3815_/A _3815_/B vssd1 vssd1 vccd1 vccd1 _3816_/A sky130_fd_sc_hd__or2_1
X_4794_ _4794_/A _4829_/A vssd1 vssd1 vccd1 vccd1 _4802_/B sky130_fd_sc_hd__and2_1
X_3745_ _3746_/A _3746_/B vssd1 vssd1 vccd1 vccd1 _3747_/A sky130_fd_sc_hd__nor2_1
X_6533_ _6533_/A _3243_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_20_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _4019_/A vssd1 vssd1 vccd1 vccd1 _3940_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5415_ _5412_/A _5412_/B _5414_/Y vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__3255__A _3257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6294__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5346_ _5541_/B _5346_/B vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__xnor2_4
X_5277_ _5277_/A _5277_/B vssd1 vssd1 vccd1 vccd1 _5300_/A sky130_fd_sc_hd__xnor2_2
XFILLER_102_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4228_ _5320_/A _4337_/B _4337_/C vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__and3_1
XFILLER_75_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ _4167_/A _4167_/B vssd1 vssd1 vccd1 vccd1 _4168_/C sky130_fd_sc_hd__xor2_4
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6560__76 vssd1 vssd1 vccd1 vccd1 _6560__76/HI _6560_/A sky130_fd_sc_hd__conb_1
XFILLER_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5975__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3530_ _6285_/Q vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3461_ _3483_/B _4814_/B _3400_/X vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__o21a_1
X_5200_ _5215_/C _5200_/B vssd1 vssd1 vccd1 vccd1 _5242_/A sky130_fd_sc_hd__xnor2_2
X_6180_ _6180_/A vssd1 vssd1 vccd1 vccd1 _6349_/D sky130_fd_sc_hd__clkbuf_1
X_3392_ _5685_/A vssd1 vssd1 vccd1 vccd1 _5701_/B sky130_fd_sc_hd__inv_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5131_ _5091_/Y _5129_/Y _5130_/X vssd1 vssd1 vccd1 vccd1 _5159_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5062_ _5062_/A _5075_/A vssd1 vssd1 vccd1 vccd1 _5114_/B sky130_fd_sc_hd__or2b_1
XFILLER_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ _4018_/A _4018_/B vssd1 vssd1 vccd1 vccd1 _4016_/B sky130_fd_sc_hd__or2_1
XFILLER_84_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4337__C _4337_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5964_ _3379_/A _5963_/X _5952_/X vssd1 vssd1 vccd1 vccd1 _5964_/Y sky130_fd_sc_hd__a21oi_1
X_4915_ _5087_/A _5087_/B _4914_/X vssd1 vssd1 vccd1 vccd1 _5066_/B sky130_fd_sc_hd__a21o_1
X_5895_ _5895_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5895_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4777_ _4805_/A _4805_/B _4776_/X vssd1 vssd1 vccd1 vccd1 _4778_/B sky130_fd_sc_hd__o21ba_2
XANTENNA__5465__A _6278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6516_ _6516_/A _3223_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_3728_ _5085_/A vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3659_ _3659_/A _3659_/B _3659_/C vssd1 vssd1 vccd1 vccd1 _3686_/A sky130_fd_sc_hd__nand3_1
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6378_ _6383_/CLK _6378_/D vssd1 vssd1 vccd1 vccd1 _6378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5329_ _5329_/A _5329_/B vssd1 vssd1 vccd1 vccd1 _5330_/C sky130_fd_sc_hd__xor2_1
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4700_ _4701_/B _4701_/C _4701_/A vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__o21a_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5727_/A vssd1 vssd1 vccd1 vccd1 _5680_/Y sky130_fd_sc_hd__inv_2
X_4631_ _4864_/D vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _5627_/A _4564_/B _4561_/X vssd1 vssd1 vccd1 vccd1 _4562_/Y sky130_fd_sc_hd__a21oi_1
X_4493_ _4493_/A _4493_/B vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__xor2_4
X_3513_ _3513_/A _3513_/B vssd1 vssd1 vccd1 vccd1 _3640_/B sky130_fd_sc_hd__xor2_1
X_6524__43 vssd1 vssd1 vccd1 vccd1 _6524__43/HI _6524_/A sky130_fd_sc_hd__conb_1
X_6301_ _6335_/CLK _6301_/D vssd1 vssd1 vccd1 vccd1 _6301_/Q sky130_fd_sc_hd__dfxtp_1
X_6232_ _6232_/A _6254_/B vssd1 vssd1 vccd1 vccd1 _6368_/D sky130_fd_sc_hd__nor2_1
X_3444_ _3556_/B vssd1 vssd1 vccd1 vccd1 _4877_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4629__A _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375_ _4815_/A vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6187_/A input7/X vssd1 vssd1 vccd1 vccd1 _6164_/A sky130_fd_sc_hd__and2_1
XFILLER_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5114_ _5114_/A _5114_/B _5114_/C vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__and3_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6094_ _6315_/Q _6189_/B vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__and2_1
XFILLER_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5045_ _5047_/A _5047_/B vssd1 vssd1 vccd1 vccd1 _5056_/B sky130_fd_sc_hd__and2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _5957_/B vssd1 vssd1 vccd1 vccd1 _5966_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5878_ _5741_/A _5891_/B _5866_/X vssd1 vssd1 vccd1 vccd1 _5879_/B sky130_fd_sc_hd__a21oi_1
X_4829_ _4829_/A _4829_/B _4852_/C vssd1 vssd1 vccd1 vccd1 _4833_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4390__A2 _4370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4539__A _5724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3443__A _6291_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4168__B _4168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5271__C _5444_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5801_ _5801_/A _6368_/Q _5801_/C vssd1 vssd1 vccd1 vccd1 _5801_/X sky130_fd_sc_hd__or3_1
XFILLER_50_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3993_ _3993_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5732_ _5732_/A _5732_/B vssd1 vssd1 vccd1 vccd1 _5732_/Y sky130_fd_sc_hd__nor2_1
X_5663_ _5618_/A _5618_/B _5626_/X _5662_/X vssd1 vssd1 vccd1 vccd1 _5663_/X sky130_fd_sc_hd__a2bb2o_1
X_4614_ _4605_/A _4613_/X _4612_/A _4612_/B _4605_/B vssd1 vssd1 vccd1 vccd1 _4614_/X
+ sky130_fd_sc_hd__a2111o_1
X_5594_ _5669_/A _5669_/B _5601_/A _5593_/X vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__a2bb2o_1
X_4545_ _4545_/A _4545_/B vssd1 vssd1 vccd1 vccd1 _4546_/C sky130_fd_sc_hd__xor2_1
XFILLER_116_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476_ _4066_/A _4067_/X _4016_/B _4018_/Y vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__o211a_1
XANTENNA__3263__A _3263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6215_ _6254_/B _6215_/B _6221_/C vssd1 vssd1 vccd1 vccd1 _6362_/D sky130_fd_sc_hd__nor3_1
X_3427_ _6301_/Q vssd1 vssd1 vccd1 vccd1 _6040_/A sky130_fd_sc_hd__buf_2
X_3358_ _3696_/A vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__clkbuf_2
X_6146_ _6335_/Q _6146_/B vssd1 vssd1 vccd1 vccd1 _6147_/A sky130_fd_sc_hd__and2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3294_/A sky130_fd_sc_hd__buf_8
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6077_ _6077_/A vssd1 vssd1 vccd1 vccd1 _6310_/D sky130_fd_sc_hd__clkbuf_1
X_5028_ _5028_/A _5028_/B vssd1 vssd1 vccd1 vccd1 _5042_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4363__A2 _4153_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _5410_/A _4301_/B _4361_/B _5440_/A vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4261_ _4261_/A _4261_/B vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3212_ _3214_/A vssd1 vssd1 vccd1 vccd1 _3212_/Y sky130_fd_sc_hd__inv_2
X_6000_ _6000_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _6001_/B sky130_fd_sc_hd__or2_1
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4192_ _3614_/B _4191_/X _3633_/X vssd1 vssd1 vccd1 vccd1 _4361_/B sky130_fd_sc_hd__a21boi_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4626__B _5710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3976_ _3976_/A _3976_/B _3976_/C vssd1 vssd1 vccd1 vccd1 _4337_/C sky130_fd_sc_hd__nand3_2
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5715_ _5715_/A _5715_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__nor2_2
X_5646_ _5646_/A _5646_/B vssd1 vssd1 vccd1 vccd1 _5646_/Y sky130_fd_sc_hd__xnor2_1
X_5577_ _5575_/A _5575_/B _5544_/X vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__a21oi_2
X_4528_ _4619_/B _4526_/Y _4619_/A vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__a21o_1
X_4459_ _4459_/A _4459_/B vssd1 vssd1 vccd1 vccd1 _4459_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6129_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6146_/B sky130_fd_sc_hd__clkbuf_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4552__A _5619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_274 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _3851_/A _3851_/B _3828_/X _3829_/X vssd1 vssd1 vccd1 vccd1 _4051_/B sky130_fd_sc_hd__a211oi_4
XFILLER_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3761_ _3807_/C _3738_/B vssd1 vssd1 vccd1 vccd1 _3805_/A sky130_fd_sc_hd__or2b_1
XFILLER_20_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6566__82 vssd1 vssd1 vccd1 vccd1 _6566__82/HI _6566_/A sky130_fd_sc_hd__conb_1
X_5500_ _5500_/A _5529_/A vssd1 vssd1 vccd1 vccd1 _5614_/A sky130_fd_sc_hd__xor2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3692_ _4714_/A _3692_/B vssd1 vssd1 vccd1 vccd1 _3734_/C sky130_fd_sc_hd__and2_2
XFILLER_9_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5431_ _5431_/A _5432_/A vssd1 vssd1 vccd1 vccd1 _5435_/B sky130_fd_sc_hd__xnor2_2
X_5362_ _5362_/A _5362_/B vssd1 vssd1 vccd1 vccd1 _5390_/A sky130_fd_sc_hd__xnor2_1
X_4313_ _5394_/A _4409_/B _5394_/B vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__and3_1
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5293_ _5294_/A _5485_/B _5505_/B _4194_/A vssd1 vssd1 vccd1 vccd1 _5322_/B sky130_fd_sc_hd__a22oi_2
X_4244_ _4388_/B vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4175_ _4177_/B _4177_/A vssd1 vssd1 vccd1 vccd1 _4175_/X sky130_fd_sc_hd__and2b_1
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _3960_/B _3960_/A vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__and2b_1
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5629_ _5629_/A _5629_/B vssd1 vssd1 vccd1 vccd1 _5630_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__B _5134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5841__A _5885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_583 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _6341_/Q _5980_/B vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__and2_1
X_4931_ _4931_/A vssd1 vssd1 vccd1 vccd1 _4933_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_439 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4862_ _4860_/A _4858_/Y _4856_/X _4857_/X vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5288__A _5486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3813_ _3813_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _3815_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3500__B1_N _3476_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _4794_/A _4793_/B _4793_/C vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__nand3_1
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3744_ _3758_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3746_/B sky130_fd_sc_hd__xnor2_1
X_6532_ _6532_/A _3242_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_3675_ _3718_/A _3718_/B vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3536__A _3536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5414_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5414_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5345_ _5345_/A _5345_/B vssd1 vssd1 vccd1 vccd1 _5346_/B sky130_fd_sc_hd__nor2_2
X_5276_ _5276_/A _5316_/B vssd1 vssd1 vccd1 vccd1 _5277_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4227_ _4227_/A _4227_/B vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__xor2_2
X_4158_ _5230_/A _4323_/B vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__nand2_2
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _4089_/A _4089_/B vssd1 vssd1 vccd1 vccd1 _4089_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4814__B _4814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4830__A _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_680 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3356__A _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3460_ _3520_/B _3548_/A _3492_/A vssd1 vssd1 vccd1 vccd1 _3463_/A sky130_fd_sc_hd__and3_1
X_3391_ _3391_/A vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__buf_2
XFILLER_97_634 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5130_ _5130_/A _5130_/B _5243_/B vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__and3_1
XFILLER_35_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5061_ _5062_/A _5061_/B _3950_/A _5038_/B vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__or4bb_1
X_4012_ _4012_/A _4012_/B vssd1 vssd1 vccd1 vccd1 _4018_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5963_ _5949_/X _5959_/X _5962_/Y _5951_/A vssd1 vssd1 vccd1 vccd1 _5963_/X sky130_fd_sc_hd__o211a_1
X_4914_ _4861_/A _4914_/B vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__and2b_1
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5894_ _5715_/A _5891_/B _5893_/Y vssd1 vssd1 vccd1 vccd1 _5895_/B sky130_fd_sc_hd__o21bai_1
X_4845_ _4844_/A _4844_/B _4866_/B vssd1 vssd1 vccd1 vccd1 _4868_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4776_ _4775_/A _4776_/B vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3727_ _5158_/A vssd1 vssd1 vccd1 vccd1 _5085_/A sky130_fd_sc_hd__clkbuf_2
X_6515_ _6515_/A _3222_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_20_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3266__A _3270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ _3657_/A _3657_/B _3657_/C vssd1 vssd1 vccd1 vccd1 _3659_/C sky130_fd_sc_hd__a21o_1
X_6377_ _6383_/CLK _6377_/D vssd1 vssd1 vccd1 vccd1 _6377_/Q sky130_fd_sc_hd__dfxtp_1
X_3589_ _4707_/A _3601_/B _3477_/D vssd1 vssd1 vccd1 vccd1 _3589_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5328_ _5328_/A _5484_/C vssd1 vssd1 vccd1 vccd1 _5329_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5259_ _5259_/A _5259_/B vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__or2_1
XFILLER_102_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4263__C _4365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4560__A _4560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_656 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4749_/A vssd1 vssd1 vccd1 vccd1 _4864_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _4560_/A _4561_/B vssd1 vssd1 vccd1 vccd1 _4561_/X sky130_fd_sc_hd__and2b_1
XFILLER_8_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6300_ _6335_/CLK _6300_/D vssd1 vssd1 vccd1 vccd1 _6300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4492_ _4492_/A _4492_/B vssd1 vssd1 vccd1 vccd1 _4493_/B sky130_fd_sc_hd__nand2_1
X_3512_ _3512_/A _3512_/B vssd1 vssd1 vccd1 vccd1 _3513_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6231_ _6367_/Q _6228_/B _6230_/Y vssd1 vssd1 vccd1 vccd1 _6367_/D sky130_fd_sc_hd__o21a_1
X_3443_ _6291_/Q _3652_/B _3652_/C _3477_/D vssd1 vssd1 vccd1 vccd1 _3446_/C sky130_fd_sc_hd__nand4_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _5904_/X _6157_/X _6158_/X _6161_/X vssd1 vssd1 vccd1 vccd1 _6341_/D sky130_fd_sc_hd__a31o_1
X_5113_ _5113_/A _5113_/B _5113_/C vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__or3_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3494_/A vssd1 vssd1 vccd1 vccd1 _4815_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _6093_/A vssd1 vssd1 vccd1 vccd1 _6315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5044_ _5042_/A _5042_/B _5078_/A vssd1 vssd1 vccd1 vccd1 _5047_/B sky130_fd_sc_hd__a21o_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5808__A1_N _5755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5946_ _5940_/A _5930_/X _5944_/Y _5945_/X vssd1 vssd1 vccd1 vccd1 _6286_/D sky130_fd_sc_hd__o211a_1
X_5877_ _5877_/A vssd1 vssd1 vccd1 vccd1 _5891_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4828_ _4840_/A _4840_/B _4840_/C vssd1 vssd1 vccd1 vccd1 _4852_/C sky130_fd_sc_hd__a21o_1
XANTENNA__5195__B _5273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4759_ _4796_/A _4820_/B _4796_/D _3601_/A vssd1 vssd1 vccd1 vccd1 _4797_/A sky130_fd_sc_hd__a22oi_4
XFILLER_108_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6584__100 vssd1 vssd1 vccd1 vccd1 _6584__100/HI _6584_/A sky130_fd_sc_hd__conb_1
XFILLER_88_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4539__B _4583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4555__A _4555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5094__A1 _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4184__B _4367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _4007_/A _4007_/B _4007_/C vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__o21ai_1
X_5800_ _6232_/A _5801_/C _5801_/A vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5731_ _5732_/A _5732_/B _6363_/Q vssd1 vssd1 vccd1 vccd1 _5731_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_50_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5662_ _5626_/A _5626_/B _5633_/X _5661_/X vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__a22o_1
X_4613_ _4613_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__or2_1
X_5593_ _5669_/A _5593_/B vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__or2_1
X_4544_ _4544_/A _4544_/B vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__xor2_1
XFILLER_116_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _4501_/A _4509_/A _4502_/B _4474_/X vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__o31ai_4
XFILLER_104_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6214_ _6362_/Q _6214_/B _6214_/C vssd1 vssd1 vccd1 vccd1 _6221_/C sky130_fd_sc_hd__and3_1
X_3426_ _3653_/B _4768_/C _4796_/D vssd1 vssd1 vccd1 vccd1 _3503_/A sky130_fd_sc_hd__o21ai_2
X_6145_ _6145_/A vssd1 vssd1 vccd1 vccd1 _6335_/D sky130_fd_sc_hd__clkbuf_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _6291_/Q vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6076_ _6309_/Q _6096_/B vssd1 vssd1 vccd1 vccd1 _6077_/A sky130_fd_sc_hd__and2_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _3903_/A _5013_/B _5013_/C vssd1 vssd1 vccd1 vccd1 _5028_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3288_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3288_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5918__B _5980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5929_ _5929_/A vssd1 vssd1 vccd1 vccd1 _5951_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4899__A1 _4726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4260_ _4260_/A _4260_/B vssd1 vssd1 vccd1 vccd1 _4467_/A sky130_fd_sc_hd__xnor2_4
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4191_ _3633_/A _3613_/B _3632_/X vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__o21ba_1
X_3211_ _3214_/A vssd1 vssd1 vccd1 vccd1 _3211_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3865__A2 _4138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _3975_/A vssd1 vssd1 vccd1 vccd1 _4337_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5714_ _5714_/A vssd1 vssd1 vccd1 vccd1 _5715_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5645_ _5875_/A _5646_/B _5644_/Y vssd1 vssd1 vccd1 vccd1 _5659_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5576_ _5683_/A _5624_/A vssd1 vssd1 vccd1 vccd1 _5576_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3274__A _3276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4527_ _4560_/A _4626_/A vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ _4553_/A _4559_/A _4457_/X vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__o21bai_1
X_3409_ _6296_/Q vssd1 vssd1 vccd1 vccd1 _6000_/A sky130_fd_sc_hd__clkbuf_2
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _4430_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6128_ _6128_/A vssd1 vssd1 vccd1 vccd1 _6329_/D sky130_fd_sc_hd__clkbuf_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__B1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6059_ _6270_/A vssd1 vssd1 vccd1 vccd1 _6254_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3760_ _3693_/A _3734_/C _3743_/B _3759_/X vssd1 vssd1 vccd1 vccd1 _3804_/A sky130_fd_sc_hd__a31o_1
XFILLER_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3691_ _3377_/A _3807_/B _3762_/B _4714_/A vssd1 vssd1 vccd1 vccd1 _3691_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5430_ _5429_/A _5449_/A _5449_/B _5448_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5432_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6581__97 vssd1 vssd1 vccd1 vccd1 _6581__97/HI _6581_/A sky130_fd_sc_hd__conb_1
XFILLER_114_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5361_ _5361_/A _5348_/X vssd1 vssd1 vccd1 vccd1 _5362_/A sky130_fd_sc_hd__or2b_1
XANTENNA__3535__A1 _3536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _4312_/A _6280_/Q _5450_/C vssd1 vssd1 vccd1 vccd1 _5394_/B sky130_fd_sc_hd__and3_1
X_5292_ _5440_/B vssd1 vssd1 vccd1 vccd1 _5505_/B sky130_fd_sc_hd__clkbuf_2
X_4243_ _3632_/X _4242_/Y _3613_/B vssd1 vssd1 vccd1 vccd1 _4388_/B sky130_fd_sc_hd__o21bai_2
X_4174_ _4165_/X _4217_/B _4173_/X vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__o21ai_1
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__A _5966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3269__A _3270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3958_ _3991_/A _3991_/B _3957_/X vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__a21bo_1
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3889_ _3902_/A _3902_/B vssd1 vssd1 vccd1 vccd1 _3905_/C sky130_fd_sc_hd__xor2_1
X_5628_ _5525_/B _5628_/B vssd1 vssd1 vccd1 vccd1 _5629_/B sky130_fd_sc_hd__and2b_1
X_5559_ _5559_/A _5559_/B vssd1 vssd1 vccd1 vccd1 _5703_/A sky130_fd_sc_hd__xor2_2
XFILLER_105_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4563__A _5619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4535__B_N _4603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _4930_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ _4861_/A _4914_/B vssd1 vssd1 vccd1 vccd1 _5087_/A sky130_fd_sc_hd__xnor2_1
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _5957_/A _3734_/B _3734_/C _3774_/B _3773_/A vssd1 vssd1 vccd1 vccd1 _3813_/B
+ sky130_fd_sc_hd__a41o_1
X_4792_ _4786_/A _4786_/B _4827_/A vssd1 vssd1 vccd1 vccd1 _4793_/C sky130_fd_sc_hd__a21o_1
X_3743_ _3743_/A _3743_/B vssd1 vssd1 vccd1 vccd1 _3758_/B sky130_fd_sc_hd__xnor2_1
X_6531_ _6531_/A _3241_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
X_3674_ _3674_/A _3674_/B vssd1 vssd1 vccd1 vccd1 _3718_/B sky130_fd_sc_hd__xnor2_2
XFILLER_9_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3536__B _3536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5413_ _6276_/Q _5469_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__and3_1
X_5344_ _5347_/A _5347_/B vssd1 vssd1 vccd1 vccd1 _5345_/B sky130_fd_sc_hd__and2b_1
XFILLER_114_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5275_ _5284_/B _5285_/B _5284_/A vssd1 vssd1 vccd1 vccd1 _5277_/A sky130_fd_sc_hd__o21ba_1
X_4226_ _4227_/A _4227_/B vssd1 vssd1 vccd1 vccd1 _4226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4367__B _4367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4157_ _4162_/B _4162_/A vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4088_ _5236_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4814__C _4814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6013__A _6187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6551__67 vssd1 vssd1 vccd1 vccd1 _6551__67/HI _6551_/A sky130_fd_sc_hd__conb_1
X_3390_ _6303_/Q vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _5059_/A _5218_/D _5059_/C vssd1 vssd1 vccd1 vccd1 _5061_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3372__A _4698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4011_ _4012_/A _4012_/B vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3426__B1 _4796_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5962_ _5957_/A _5959_/C _5949_/X vssd1 vssd1 vccd1 vccd1 _5962_/Y sky130_fd_sc_hd__o21ai_1
X_4913_ _5125_/B _5125_/C _5125_/A vssd1 vssd1 vccd1 vccd1 _5087_/B sky130_fd_sc_hd__a21bo_1
X_5893_ _5714_/A _5891_/B _5886_/A vssd1 vssd1 vccd1 vccd1 _5893_/Y sky130_fd_sc_hd__a21oi_1
X_4844_ _4844_/A _4844_/B _4866_/B vssd1 vssd1 vccd1 vccd1 _4868_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4775_ _4775_/A _4776_/B vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__xor2_2
XFILLER_21_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3726_ _4115_/A vssd1 vssd1 vccd1 vccd1 _5158_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6514_ _6514_/A _3220_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_3657_ _3657_/A _3657_/B _3657_/C vssd1 vssd1 vccd1 vccd1 _3659_/B sky130_fd_sc_hd__nand3_1
X_6376_ _6383_/CLK _6376_/D vssd1 vssd1 vccd1 vccd1 _6376_/Q sky130_fd_sc_hd__dfxtp_1
X_3588_ _3585_/B _3585_/C _3594_/B vssd1 vssd1 vccd1 vccd1 _3617_/B sky130_fd_sc_hd__o21ai_1
X_5327_ _5439_/B vssd1 vssd1 vccd1 vccd1 _5484_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3282__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _5301_/A _5301_/B vssd1 vssd1 vccd1 vccd1 _5259_/B sky130_fd_sc_hd__nor2_1
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _4167_/B _4227_/A _4187_/A _4187_/B vssd1 vssd1 vccd1 vccd1 _4210_/C sky130_fd_sc_hd__o22ai_1
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5189_ _5186_/A _5186_/Y _5148_/X _5188_/X vssd1 vssd1 vccd1 vccd1 _5189_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5672__A _5672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5893__A1 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3192__A _3195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5645__A1 _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_484 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4560_ _4560_/A _4561_/B vssd1 vssd1 vccd1 vccd1 _4564_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4491_ _4491_/A _3937_/B vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__or2b_2
X_3511_ _3508_/Y _3509_/X _3536_/A _3475_/Y vssd1 vssd1 vccd1 vccd1 _3512_/B sky130_fd_sc_hd__o211a_1
XFILLER_116_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6230_ _6367_/Q _6228_/B _5952_/X vssd1 vssd1 vccd1 vccd1 _6230_/Y sky130_fd_sc_hd__a21oi_1
X_3442_ _6287_/Q _3556_/B vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__and2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _6335_/Q _6159_/X _6160_/X _6293_/D vssd1 vssd1 vccd1 vccd1 _6161_/X sky130_fd_sc_hd__o31a_1
X_3373_ _6288_/Q vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5112_ _5107_/A _5107_/B _5107_/C vssd1 vssd1 vccd1 vccd1 _5113_/C sky130_fd_sc_hd__a21oi_1
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6140_/A input4/X vssd1 vssd1 vccd1 vccd1 _6093_/A sky130_fd_sc_hd__and2_1
XFILLER_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5043_ _5046_/B _5043_/B _5043_/C vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__and3_1
XFILLER_78_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5650__B1_N _4138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5945_ _6187_/A vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5876_ _5876_/A _5876_/B vssd1 vssd1 vccd1 vccd1 _5879_/A sky130_fd_sc_hd__nand2_1
X_4827_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4840_/C sky130_fd_sc_hd__nand2_1
X_4758_ _4758_/A _4758_/B vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4689_ _4689_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__or2b_1
X_3709_ _3730_/A _3707_/Y _3687_/Y _3688_/X vssd1 vssd1 vccd1 vccd1 _3710_/B sky130_fd_sc_hd__o211a_1
X_6515__34 vssd1 vssd1 vccd1 vccd1 _6515__34/HI _6515_/A sky130_fd_sc_hd__conb_1
XFILLER_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6359_ _6359_/CLK _6359_/D vssd1 vssd1 vccd1 vccd1 _6359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4465__B _4465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _3991_/A _3991_/B vssd1 vssd1 vccd1 vccd1 _4007_/C sky130_fd_sc_hd__xor2_1
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5730_ _3383_/A _5728_/X _5700_/X _5875_/A _5729_/Y vssd1 vssd1 vccd1 vccd1 _5732_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3468__B1_N _4818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5661_ _5633_/A _5633_/B _5639_/X _5660_/X vssd1 vssd1 vccd1 vccd1 _5661_/X sky130_fd_sc_hd__a22o_1
X_4612_ _4612_/A _4612_/B _4612_/C vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__or3_1
X_5592_ _5679_/A _5637_/A vssd1 vssd1 vccd1 vccd1 _5593_/B sky130_fd_sc_hd__and2_1
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4543_ _4543_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4612_/A sky130_fd_sc_hd__xnor2_1
X_4474_ _4141_/B _4141_/C _4141_/A vssd1 vssd1 vccd1 vccd1 _4474_/X sky130_fd_sc_hd__a21o_1
X_6213_ _6214_/B _6214_/C _6362_/Q vssd1 vssd1 vccd1 vccd1 _6215_/B sky130_fd_sc_hd__a21oi_1
X_3425_ _3387_/A _5685_/A _6301_/Q vssd1 vssd1 vccd1 vccd1 _4796_/D sky130_fd_sc_hd__a21o_2
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6144_ _6334_/Q _6146_/B vssd1 vssd1 vccd1 vccd1 _6145_/A sky130_fd_sc_hd__and2_1
X_3356_ _5955_/A _5940_/A vssd1 vssd1 vccd1 vccd1 _5691_/C sky130_fd_sc_hd__or2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6075_ _6098_/A vssd1 vssd1 vccd1 vccd1 _6096_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A _5026_/B vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__xor2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4596__A1 _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _5924_/X _5925_/Y _5926_/X _5927_/X vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__o22a_1
X_5859_ _5980_/B vssd1 vssd1 vccd1 vccd1 _6189_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _5324_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__nand2_1
X_3210_ _3214_/A vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3380__A _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4578__A1 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _5130_/A _4268_/B vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__nand2_1
X_5713_ _5890_/A _5700_/X _5712_/X _3384_/A vssd1 vssd1 vccd1 vccd1 _5713_/Y sky130_fd_sc_hd__a22oi_2
X_5644_ _5644_/A _5644_/B vssd1 vssd1 vccd1 vccd1 _5644_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5575_ _5575_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _5624_/A sky130_fd_sc_hd__xor2_4
X_4526_ _4615_/A _4615_/B vssd1 vssd1 vccd1 vccd1 _4526_/Y sky130_fd_sc_hd__nand2_1
X_4457_ _4425_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4457_/X sky130_fd_sc_hd__and2b_1
X_3408_ _3405_/X _3406_/X _6295_/Q _3517_/A vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__a211oi_2
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input7_A io_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4388_ _5440_/A _4388_/B _5484_/B vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__and3_1
X_6127_ _6328_/Q _6127_/B vssd1 vssd1 vccd1 vccd1 _6128_/A sky130_fd_sc_hd__and2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3290__A _3294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _6285_/Q vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6058_ _6061_/A _6023_/X _6055_/X _6057_/Y _5904_/X vssd1 vssd1 vccd1 vccd1 _6303_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5172_/B vssd1 vssd1 vccd1 vccd1 _5316_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3449__B _4814_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5945__A _6187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_192 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6016__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _3690_/A vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5360_ _5360_/A _5360_/B vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3535__A2 _3536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4311_ _4311_/A _4311_/B vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__nor2_1
X_5291_ _5291_/A vssd1 vssd1 vccd1 vccd1 _5440_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4242_ _3632_/A _3632_/C _5325_/C vssd1 vssd1 vccd1 vccd1 _4242_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _4216_/A _4216_/B vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__or2b_1
XFILLER_95_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4934__A _5966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _3957_/A _3949_/B vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__or2b_1
X_6557__73 vssd1 vssd1 vccd1 vccd1 _6557__73/HI _6557_/A sky130_fd_sc_hd__conb_1
X_3888_ _4925_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _3902_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3285__A _3288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5627_ _5627_/A _5627_/B vssd1 vssd1 vccd1 vccd1 _5633_/A sky130_fd_sc_hd__xnor2_1
X_5558_ _5560_/B _5561_/B _5560_/A vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__o21bai_4
X_4509_ _4509_/A _4509_/B vssd1 vssd1 vccd1 vccd1 _4510_/B sky130_fd_sc_hd__nor2_2
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5489_ _5489_/A _5489_/B vssd1 vssd1 vccd1 vccd1 _5490_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6312__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3907__B _4138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3195__A _3195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4860_/A _4860_/B vssd1 vssd1 vccd1 vccd1 _4914_/B sky130_fd_sc_hd__or2_1
X_3811_ _3811_/A _3811_/B vssd1 vssd1 vccd1 vccd1 _3813_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6530_ _6530_/A _3239_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
X_4791_ _4791_/A _4791_/B vssd1 vssd1 vccd1 vccd1 _4793_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3756__A2 _4168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3742_ _3759_/B _3742_/B vssd1 vssd1 vccd1 vccd1 _3743_/B sky130_fd_sc_hd__xnor2_1
XFILLER_9_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3673_ _3673_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3674_/B sky130_fd_sc_hd__nor2_1
X_5412_ _5412_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__xor2_1
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5343_ _5343_/A _5343_/B vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__xnor2_2
XFILLER_114_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5274_ _5274_/A _5312_/A _5274_/C _5274_/D vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__and4_1
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6335__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4225_ _5274_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4227_/B sky130_fd_sc_hd__nand2_2
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4162_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _4095_/A _4095_/B vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4989_ _4989_/A _4989_/B vssd1 vssd1 vccd1 vccd1 _5024_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_410 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4935__A1 _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6358__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4010_ _4010_/A _4010_/B vssd1 vssd1 vccd1 vccd1 _4012_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_330 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5961_ _5957_/A _5930_/X _5960_/Y _5945_/X vssd1 vssd1 vccd1 vccd1 _6288_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4912_ _4873_/A _4910_/A _4860_/B _4862_/X vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__a211o_1
XFILLER_21_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5892_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__nor2_1
X_4843_ _4877_/A _4877_/C vssd1 vssd1 vccd1 vccd1 _4866_/B sky130_fd_sc_hd__nand2_1
X_4774_ _4783_/A _4783_/B _4773_/X vssd1 vssd1 vccd1 vccd1 _4776_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3725_ _5246_/A vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6513_ _6513_/A _3219_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
X_3656_ _3688_/A _3688_/B vssd1 vssd1 vccd1 vccd1 _3657_/C sky130_fd_sc_hd__xor2_1
X_6375_ _6375_/CLK _6375_/D vssd1 vssd1 vccd1 vccd1 _6375_/Q sky130_fd_sc_hd__dfxtp_1
X_3587_ _3619_/A _3619_/B vssd1 vssd1 vccd1 vccd1 _3626_/A sky130_fd_sc_hd__xor2_2
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _4312_/A _3632_/C _5289_/A _5325_/X vssd1 vssd1 vccd1 vccd1 _5439_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_6__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5257_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5301_/B sky130_fd_sc_hd__xor2_1
XFILLER_102_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4208_ _5312_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4227_/A sky130_fd_sc_hd__nand2_2
XFILLER_87_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5188_ _5151_/B _5148_/C _5187_/Y _5141_/X vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4139_ _4139_/A _4139_/B vssd1 vssd1 vccd1 vccd1 _4142_/C sky130_fd_sc_hd__xnor2_1
XFILLER_56_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5342__A1 _4062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__A _4569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3510_ _3536_/A _3475_/Y _3508_/Y _3509_/X vssd1 vssd1 vccd1 vccd1 _3512_/A sky130_fd_sc_hd__a211oi_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4490_ _4490_/A _4490_/B vssd1 vssd1 vccd1 vccd1 _5702_/A sky130_fd_sc_hd__xnor2_4
XFILLER_7_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3441_ _3547_/B vssd1 vssd1 vccd1 vccd1 _3556_/B sky130_fd_sc_hd__clkbuf_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _6338_/Q _6337_/Q _6340_/Q _6339_/Q vssd1 vssd1 vccd1 vccd1 _6160_/X sky130_fd_sc_hd__or4_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3372_ _4698_/A vssd1 vssd1 vccd1 vccd1 _3379_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5111_ _5118_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__or2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _5861_/X _6084_/X _6085_/X _6088_/X _6384_/D vssd1 vssd1 vccd1 vccd1 _6314_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5042_ _5042_/A _5042_/B vssd1 vssd1 vccd1 vccd1 _5043_/C sky130_fd_sc_hd__xor2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5970_/A _5944_/B vssd1 vssd1 vccd1 vccd1 _5944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5875_ _5875_/A _5877_/A vssd1 vssd1 vccd1 vccd1 _5876_/B sky130_fd_sc_hd__or2_1
X_4826_ _4785_/A _4785_/C _4768_/D _3601_/A vssd1 vssd1 vccd1 vccd1 _4827_/B sky130_fd_sc_hd__a22o_1
XANTENNA__3558__A _4865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4757_/A _4757_/B _4757_/C vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__and3_1
X_4688_ _4742_/A _4742_/B vssd1 vssd1 vccd1 vccd1 _4743_/A sky130_fd_sc_hd__or2_1
X_3708_ _3687_/Y _3688_/X _3730_/A _3707_/Y vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__a211oi_1
XFILLER_4_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3639_ _3941_/A _3975_/A vssd1 vssd1 vccd1 vccd1 _3718_/A sky130_fd_sc_hd__nor2b_2
XANTENNA__3293__A _3294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6530__49 vssd1 vssd1 vccd1 vccd1 _6530__49/HI _6530_/A sky130_fd_sc_hd__conb_1
X_6358_ _6384_/CLK _6358_/D vssd1 vssd1 vccd1 vccd1 _6358_/Q sky130_fd_sc_hd__dfxtp_1
X_5309_ _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5310_/B sky130_fd_sc_hd__xnor2_2
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_49 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_444 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6289_ _6335_/CLK _6289_/D vssd1 vssd1 vccd1 vccd1 _6289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_48 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _4040_/A _4040_/B vssd1 vssd1 vccd1 vccd1 _4007_/B sky130_fd_sc_hd__and2_1
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5660_ _5639_/A _5639_/B _5658_/Y _5659_/Y vssd1 vssd1 vccd1 vccd1 _5660_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4611_ _4611_/A _4611_/B _4611_/C _4611_/D vssd1 vssd1 vccd1 vccd1 _4612_/C sky130_fd_sc_hd__or4_1
X_5591_ _5727_/A _5644_/A vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__or2_1
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4542_ _4544_/A _4542_/B vssd1 vssd1 vccd1 vccd1 _4542_/X sky130_fd_sc_hd__or2_1
X_4473_ _4512_/A _4512_/B _4509_/B _4472_/Y vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__a211oi_4
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3424_ _4707_/B vssd1 vssd1 vccd1 vccd1 _4768_/C sky130_fd_sc_hd__clkbuf_2
X_6212_ _6214_/B _6214_/C _6211_/Y vssd1 vssd1 vccd1 vccd1 _6361_/D sky130_fd_sc_hd__o21a_1
X_6143_ _6143_/A vssd1 vssd1 vccd1 vccd1 _6334_/D sky130_fd_sc_hd__clkbuf_1
X_3355_ _4726_/A vssd1 vssd1 vccd1 vccd1 _5940_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3286_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3286_/Y sky130_fd_sc_hd__inv_2
X_6074_ _6074_/A vssd1 vssd1 vccd1 vccd1 _6309_/D sky130_fd_sc_hd__clkbuf_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__B1 _4818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _5557_/A _5557_/B vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__nor2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4672__A _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_355 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6034__A2 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5927_ _6332_/Q _6341_/Q vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3288__A _3288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5858_ input8/X vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__inv_2
X_4809_ _4812_/A _4812_/B vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__or2b_1
X_5789_ _3384_/A _5788_/X _5778_/X _5733_/X vssd1 vssd1 vccd1 vccd1 _5791_/B sky130_fd_sc_hd__a22oi_1
XFILLER_5_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3751__A _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4582__A _4583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3198__A _3201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3973_ _3973_/A vssd1 vssd1 vccd1 vccd1 _4268_/B sky130_fd_sc_hd__clkbuf_2
X_5712_ _3396_/Y _5710_/X _5711_/Y _5687_/X vssd1 vssd1 vccd1 vccd1 _5712_/X sky130_fd_sc_hd__a22o_1
X_5643_ _5644_/A _5644_/B vssd1 vssd1 vccd1 vccd1 _5646_/B sky130_fd_sc_hd__xor2_1
X_5574_ _5737_/B vssd1 vssd1 vccd1 vccd1 _5574_/Y sky130_fd_sc_hd__inv_2
X_4525_ _5710_/A _4569_/A vssd1 vssd1 vccd1 vccd1 _4615_/B sky130_fd_sc_hd__xnor2_1
X_4456_ _4558_/B _4566_/A _4558_/A vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__a21o_1
X_4387_ _5465_/B vssd1 vssd1 vccd1 vccd1 _5484_/B sky130_fd_sc_hd__clkbuf_1
X_6500__19 vssd1 vssd1 vccd1 vccd1 _6500__19/HI _6500_/A sky130_fd_sc_hd__conb_1
X_3407_ _6294_/Q vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__clkbuf_2
X_6126_ _6126_/A vssd1 vssd1 vccd1 vccd1 _6328_/D sky130_fd_sc_hd__clkbuf_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _4933_/A vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4386__B _5511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3269_ _3270_/A vssd1 vssd1 vccd1 vccd1 _3269_/Y sky130_fd_sc_hd__inv_2
X_6057_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6057_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5008_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _5172_/B sky130_fd_sc_hd__xor2_4
XFILLER_66_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4577__A _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3481__A _6291_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4310_ _5330_/A _4389_/A _4281_/C vssd1 vssd1 vccd1 vccd1 _4311_/B sky130_fd_sc_hd__a21oi_1
X_5290_ _5290_/A _5290_/B vssd1 vssd1 vccd1 vccd1 _5291_/A sky130_fd_sc_hd__or2_1
X_4241_ _5330_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__nand2_1
X_4172_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3956_ _3956_/A _3956_/B vssd1 vssd1 vccd1 vccd1 _3991_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4950__A _5966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _4929_/A _4166_/B vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__nand2_1
X_5626_ _5626_/A _5626_/B vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__or2_1
X_5557_ _5557_/A _5557_/B vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__and2_1
X_6572__88 vssd1 vssd1 vccd1 vccd1 _6572__88/HI _6572_/A sky130_fd_sc_hd__conb_1
X_4508_ _4512_/A _4512_/B _4472_/Y vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__a21oi_2
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5488_ _5488_/A _5488_/B vssd1 vssd1 vccd1 vccd1 _5490_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4439_ _4558_/B _4439_/B vssd1 vssd1 vccd1 vccd1 _4565_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6320_/Q _6319_/Q _6322_/Q _6321_/Q vssd1 vssd1 vccd1 vccd1 _6110_/C sky130_fd_sc_hd__and4_1
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5675__B _5675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5911__A1 _5906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6287__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _3810_/A _3810_/B _3810_/C vssd1 vssd1 vccd1 vccd1 _3811_/B sky130_fd_sc_hd__and3_1
XFILLER_60_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4790_ _4820_/A _4877_/C vssd1 vssd1 vccd1 vccd1 _4791_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5866__A _5866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ _3741_/A _3741_/B vssd1 vssd1 vccd1 vccd1 _3742_/B sky130_fd_sc_hd__xor2_1
XFILLER_32_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _3672_/A _3672_/B _3672_/C vssd1 vssd1 vccd1 vccd1 _3673_/B sky130_fd_sc_hd__and3_1
XFILLER_70_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5411_ _5411_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__nand2_1
X_5342_ _4062_/A _5355_/B _5315_/A _5341_/Y vssd1 vssd1 vccd1 vccd1 _5347_/A sky130_fd_sc_hd__a31oi_4
XFILLER_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _5320_/A _5273_/B vssd1 vssd1 vccd1 vccd1 _5285_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4224_ _4224_/A _4224_/B vssd1 vssd1 vccd1 vccd1 _4469_/A sky130_fd_sc_hd__xnor2_4
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4155_ _5243_/A _4367_/B _4115_/C vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__a21oi_1
XFILLER_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4945__A _5059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4086_ _4086_/A _4086_/B vssd1 vssd1 vccd1 vccd1 _4095_/B sky130_fd_sc_hd__or2_1
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5197__A2 _5358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_678 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4988_ _4988_/A _4988_/B _4988_/C vssd1 vssd1 vccd1 vccd1 _4989_/B sky130_fd_sc_hd__nor3_1
X_3939_ _3939_/A _3939_/B vssd1 vssd1 vccd1 vccd1 _3960_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3296__A _3300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5609_ _5605_/Y _5613_/B _5608_/X vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__o21a_1
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6589_ _6589_/A _3308_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4871__A1 _4865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _5958_/Y _5959_/X _5970_/A vssd1 vssd1 vccd1 vccd1 _5960_/Y sky130_fd_sc_hd__o21ai_1
X_4911_ _4892_/X _4909_/X _5161_/A vssd1 vssd1 vccd1 vccd1 _5125_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5891_ _5899_/A _5891_/B vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__nor2_1
X_4842_ _4842_/A _4842_/B _4864_/C _4864_/D vssd1 vssd1 vccd1 vccd1 _4844_/B sky130_fd_sc_hd__nand4_2
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _4772_/A _4773_/B vssd1 vssd1 vccd1 vccd1 _4773_/X sky130_fd_sc_hd__and2b_1
X_6512_ _6512_/A _3218_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
X_3724_ _5330_/A vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__buf_2
X_3655_ _4820_/A _3762_/B _3495_/B _3654_/Y vssd1 vssd1 vccd1 vccd1 _3688_/B sky130_fd_sc_hd__a31o_1
XFILLER_9_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6542__58 vssd1 vssd1 vccd1 vccd1 _6542__58/HI _6542_/A sky130_fd_sc_hd__conb_1
X_6374_ _6375_/CLK _6374_/D vssd1 vssd1 vccd1 vccd1 _6374_/Q sky130_fd_sc_hd__dfxtp_1
X_3586_ _3585_/B _3617_/A vssd1 vssd1 vccd1 vccd1 _3619_/B sky130_fd_sc_hd__and2b_1
XFILLER_114_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5325_ _5935_/A _5325_/B _5325_/C vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__or3_1
X_5256_ _5256_/A _5256_/B vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__xor2_2
X_4207_ _5278_/A _4207_/B vssd1 vssd1 vccd1 vccd1 _4213_/A sky130_fd_sc_hd__nand2_2
XFILLER_102_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5187_ _5141_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4138_ _4138_/A _4138_/B _4138_/C vssd1 vssd1 vccd1 vccd1 _4142_/B sky130_fd_sc_hd__and3_1
XANTENNA__4394__B _4412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4069_ _4531_/B vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__inv_2
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4090__A2 _3947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5342__A2 _5355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4585__A _5001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3440_ _3405_/X _6303_/Q _3517_/A vssd1 vssd1 vccd1 vccd1 _3547_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6040__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3371_ _4644_/A vssd1 vssd1 vccd1 vccd1 _4698_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5110_ _5109_/A _5145_/B _5109_/C vssd1 vssd1 vccd1 vccd1 _5111_/B sky130_fd_sc_hd__a21oi_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _6090_/A vssd1 vssd1 vccd1 vccd1 _6384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5041_ _5040_/A _5040_/B _3877_/A _5145_/B vssd1 vssd1 vccd1 vccd1 _5043_/B sky130_fd_sc_hd__a2bb2o_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5943_ _5943_/A _5943_/B vssd1 vssd1 vccd1 vccd1 _5944_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6215__A _6254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5874_ _5875_/A _5877_/A vssd1 vssd1 vccd1 vccd1 _5876_/A sky130_fd_sc_hd__nand2_1
X_4825_ _4818_/B _4816_/B _4816_/C vssd1 vssd1 vccd1 vccd1 _4840_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4756_ _4757_/A _4757_/B _4757_/C vssd1 vssd1 vccd1 vccd1 _4758_/A sky130_fd_sc_hd__a21oi_1
X_4687_ _4687_/A _4687_/B vssd1 vssd1 vccd1 vccd1 _4742_/B sky130_fd_sc_hd__xnor2_1
X_3707_ _3731_/B _3706_/C _3706_/A vssd1 vssd1 vccd1 vccd1 _3707_/Y sky130_fd_sc_hd__a21oi_1
X_3638_ _3976_/A _3976_/C _3976_/B vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__a21o_1
X_3569_ _3621_/A _3621_/B _3621_/C vssd1 vssd1 vccd1 vccd1 _3624_/B sky130_fd_sc_hd__o21ai_2
X_6357_ _6357_/CLK _6357_/D vssd1 vssd1 vccd1 vccd1 _6357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5308_ _5544_/B _5308_/B vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6288_ _6335_/CLK _6288_/D vssd1 vssd1 vccd1 vccd1 _6288_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5239_ _5221_/B _5221_/C _5221_/D _5221_/A vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__o22a_1
XFILLER_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5013__B _5013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6591__107 vssd1 vssd1 vccd1 vccd1 _6591__107/HI _6591_/A sky130_fd_sc_hd__conb_1
XFILLER_12_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3574__A1 _3601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6506__25 vssd1 vssd1 vccd1 vccd1 _6506__25/HI _6506_/A sky130_fd_sc_hd__conb_1
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4826__B2 _3601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4610_ _4550_/X _4556_/Y _4608_/X _4609_/Y vssd1 vssd1 vccd1 vccd1 _4611_/D sky130_fd_sc_hd__a211o_1
XANTENNA__5874__A _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5590_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__xnor2_2
X_4541_ _4543_/A _4543_/B _4544_/B vssd1 vssd1 vccd1 vccd1 _4542_/B sky130_fd_sc_hd__o21ba_1
X_4472_ _4472_/A _4472_/B vssd1 vssd1 vccd1 vccd1 _4472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6211_ _6214_/B _6214_/C _5952_/X vssd1 vssd1 vccd1 vccd1 _6211_/Y sky130_fd_sc_hd__a21oi_1
X_3423_ _3458_/A vssd1 vssd1 vccd1 vccd1 _3653_/B sky130_fd_sc_hd__clkbuf_2
X_6142_ _6333_/Q _6146_/B vssd1 vssd1 vccd1 vccd1 _6143_/A sky130_fd_sc_hd__and2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3661_/A vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__buf_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__inv_2
X_6073_ _6308_/Q _6073_/B vssd1 vssd1 vccd1 vccd1 _6074_/A sky130_fd_sc_hd__and2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5024_ _5024_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5557_/B sky130_fd_sc_hd__xnor2_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4672__B _4726_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5926_ _6341_/Q _6332_/Q vssd1 vssd1 vccd1 vccd1 _5926_/X sky130_fd_sc_hd__and2b_1
XFILLER_110_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5857_ _5868_/A vssd1 vssd1 vccd1 vccd1 _5857_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4808_ _4808_/A _4808_/B vssd1 vssd1 vccd1 vccd1 _4812_/B sky130_fd_sc_hd__xnor2_2
X_5788_ _5769_/X _5727_/Y _5771_/Y _5724_/Y vssd1 vssd1 vccd1 vccd1 _5788_/X sky130_fd_sc_hd__a22o_1
X_4739_ _4745_/B _4739_/B vssd1 vssd1 vccd1 vccd1 _4747_/B sky130_fd_sc_hd__or2_2
XFILLER_107_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3859__A2 _4166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578__94 vssd1 vssd1 vccd1 vccd1 _6578__94/HI _6578_/A sky130_fd_sc_hd__conb_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5588__B _5630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _3972_/A _3972_/B vssd1 vssd1 vccd1 vccd1 _3984_/A sky130_fd_sc_hd__xnor2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5711_ _5711_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5711_/Y sky130_fd_sc_hd__xnor2_1
X_5642_ _5642_/A _5642_/B vssd1 vssd1 vccd1 vccd1 _5644_/B sky130_fd_sc_hd__nand2_1
X_5573_ _5676_/A _5675_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5737_/B sky130_fd_sc_hd__or3_1
XFILLER_116_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4524_ _4624_/A _4577_/A vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__and2_1
XFILLER_116_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6497__16 vssd1 vssd1 vccd1 vccd1 _6497__16/HI _6497_/A sky130_fd_sc_hd__conb_1
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4455_ _4455_/A _4455_/B vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__xnor2_1
XFILLER_116_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4386_ _4386_/A _5511_/B vssd1 vssd1 vccd1 vccd1 _5465_/B sky130_fd_sc_hd__nor2_1
X_3406_ _6303_/Q vssd1 vssd1 vccd1 vccd1 _3406_/X sky130_fd_sc_hd__buf_2
XFILLER_98_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3337_ _4694_/A vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__clkbuf_2
X_6125_ _6327_/Q _6127_/B vssd1 vssd1 vccd1 vccd1 _6126_/A sky130_fd_sc_hd__and2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3268_ _3270_/A vssd1 vssd1 vccd1 vccd1 _3268_/Y sky130_fd_sc_hd__inv_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6055_/A _6060_/C _6055_/C vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__a21o_1
X_5007_ _5007_/A _5180_/D vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3199_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3199_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3299__A _3300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5909_ _5909_/A _5909_/B vssd1 vssd1 vccd1 vccd1 _5910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6597__113 vssd1 vssd1 vccd1 vccd1 _6597__113/HI _6597_/A sky130_fd_sc_hd__conb_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4240_ _4240_/A _4240_/B vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__nand2_1
X_4171_ _4180_/A _4170_/X vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__or2b_1
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_215 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5599__A _5737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3955_ _3993_/A _3961_/B _3954_/X vssd1 vssd1 vccd1 vccd1 _3956_/B sky130_fd_sc_hd__o21a_1
X_3886_ _5013_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _3890_/A sky130_fd_sc_hd__nand2_1
X_5625_ _5755_/A _5627_/B _5624_/X vssd1 vssd1 vccd1 vccd1 _5626_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5905__C1 _5904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5556_ _5562_/A _5562_/B _5055_/A vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__a21oi_2
X_4507_ _4621_/A _4621_/B vssd1 vssd1 vccd1 vccd1 _5735_/B sky130_fd_sc_hd__nand2_1
X_5487_ _5505_/C _5504_/A vssd1 vssd1 vccd1 vccd1 _5488_/B sky130_fd_sc_hd__nor2_1
X_4438_ _4438_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4439_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4369_ _4369_/A _4369_/B vssd1 vssd1 vccd1 vccd1 _4380_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6108_ _6108_/A vssd1 vssd1 vccd1 vccd1 _6322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6039_ _6300_/Q _6023_/X _6038_/X _6013_/X vssd1 vssd1 vccd1 vccd1 _6300_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5436__B2 _6278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_654 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3757__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6548__64 vssd1 vssd1 vccd1 vccd1 _6548__64/HI _6548_/A sky130_fd_sc_hd__conb_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4588__A _4603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5691__B _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _3740_/A _3740_/B vssd1 vssd1 vccd1 vccd1 _3741_/B sky130_fd_sc_hd__xor2_1
XFILLER_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3671_ _3672_/A _3672_/B _3672_/C vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__a21oi_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5410_ _5410_/A _5410_/B vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__nand2_1
X_5341_ _5341_/A _5341_/B vssd1 vssd1 vccd1 vccd1 _5341_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5272_ _5231_/B _5426_/B _5271_/X vssd1 vssd1 vccd1 vccd1 _5284_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4223_ _4472_/A _4472_/B vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__xor2_4
X_4154_ _4189_/A _4188_/B _4188_/A vssd1 vssd1 vccd1 vccd1 _4162_/B sky130_fd_sc_hd__o21ba_1
XFILLER_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4085_ _4052_/B _4038_/C _4038_/A vssd1 vssd1 vccd1 vccd1 _4086_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6218__A _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6091__A1 _5861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4987_ _4988_/A _4988_/B _4988_/C vssd1 vssd1 vccd1 vccd1 _4989_/A sky130_fd_sc_hd__o21a_1
X_3938_ _3938_/A _3938_/B _3938_/C vssd1 vssd1 vccd1 vccd1 _4479_/C sky130_fd_sc_hd__nand3_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3869_ _5037_/A _3906_/B vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6588_ _6588_/A _3306_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_5608_ _5675_/B _5608_/B vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__or2_1
X_5539_ _5378_/B _5539_/B vssd1 vssd1 vccd1 vccd1 _5539_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4910_ _4910_/A _4910_/B _4910_/C vssd1 vssd1 vccd1 vccd1 _5161_/A sky130_fd_sc_hd__and3_1
X_5890_ _5890_/A _5899_/B vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__and2_1
XFILLER_45_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4841_ _4842_/A _4879_/D _4864_/D _4879_/A vssd1 vssd1 vccd1 vccd1 _4844_/A sky130_fd_sc_hd__a22o_1
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772_ _4772_/A _4773_/B vssd1 vssd1 vccd1 vccd1 _4783_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6511_ _6511_/A _3217_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
X_3723_ _6279_/Q vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3654_ _3687_/A _3693_/A vssd1 vssd1 vccd1 vccd1 _3654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6373_ _6375_/CLK _6373_/D vssd1 vssd1 vccd1 vccd1 _6373_/Q sky130_fd_sc_hd__dfxtp_1
X_3585_ _3594_/B _3585_/B _3585_/C vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__or3_1
XFILLER_114_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5324_ _5324_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__nand2_1
X_5255_ _5255_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5256_/B sky130_fd_sc_hd__nand2_1
X_4206_ _4214_/B _4206_/B vssd1 vssd1 vccd1 vccd1 _4233_/A sky130_fd_sc_hd__xnor2_4
X_5186_ _5186_/A _5186_/B _5186_/C _5186_/D vssd1 vssd1 vccd1 vccd1 _5186_/Y sky130_fd_sc_hd__nand4_2
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4137_/A _4137_/B vssd1 vssd1 vccd1 vccd1 _4142_/A sky130_fd_sc_hd__and2_1
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4068_ _4016_/B _4018_/Y _4066_/A _4067_/X vssd1 vssd1 vccd1 vccd1 _4531_/B sky130_fd_sc_hd__a211oi_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_55 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4866__A _4898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3945__A _5064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3370_ _4820_/A vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5040_ _5040_/A _5040_/B _3877_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__or4bb_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5942_ _3381_/B _5957_/B _5936_/X vssd1 vssd1 vccd1 vccd1 _5943_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5873_ _5741_/A _5857_/X _5869_/Y _5872_/X vssd1 vssd1 vccd1 vccd1 _6275_/D sky130_fd_sc_hd__o211a_1
X_4824_ _4794_/A _4793_/C _4793_/B vssd1 vssd1 vccd1 vccd1 _4829_/B sky130_fd_sc_hd__a21o_1
X_4755_ _4755_/A _4755_/B vssd1 vssd1 vccd1 vccd1 _4757_/C sky130_fd_sc_hd__nor2_1
X_3706_ _3706_/A _3731_/B _3706_/C vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__and3_1
X_4686_ _4686_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__nor2_1
X_3637_ _4022_/A _4071_/A vssd1 vssd1 vccd1 vccd1 _3976_/B sky130_fd_sc_hd__or2_1
XFILLER_115_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6356_ _6357_/CLK _6356_/D vssd1 vssd1 vccd1 vccd1 _6356_/Q sky130_fd_sc_hd__dfxtp_1
X_3568_ _3570_/A _3570_/B _3567_/X vssd1 vssd1 vccd1 vccd1 _3621_/C sky130_fd_sc_hd__a21oi_1
X_5307_ _5310_/A _5305_/X _5306_/X vssd1 vssd1 vccd1 vccd1 _5308_/B sky130_fd_sc_hd__o21ba_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3499_ _3476_/Y _3642_/B _3499_/C vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__and3b_1
X_6287_ _6335_/CLK _6287_/D vssd1 vssd1 vccd1 vccd1 _6287_/Q sky130_fd_sc_hd__dfxtp_1
X_5238_ _5235_/A _5235_/B _5237_/Y vssd1 vssd1 vccd1 vccd1 _5268_/A sky130_fd_sc_hd__o21ba_2
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5169_ _5169_/A _5169_/B vssd1 vssd1 vccd1 vccd1 _5202_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4299__C _4365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _5724_/A _4583_/A vssd1 vssd1 vccd1 vccd1 _4544_/B sky130_fd_sc_hd__nor2_1
X_4471_ _4175_/X _4181_/A _4141_/C _4142_/X vssd1 vssd1 vccd1 vccd1 _4509_/B sky130_fd_sc_hd__o211a_1
XFILLER_7_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3422_ _3692_/B vssd1 vssd1 vccd1 vccd1 _3807_/B sky130_fd_sc_hd__clkbuf_2
X_6210_ _6214_/C _6254_/B vssd1 vssd1 vccd1 vccd1 _6360_/D sky130_fd_sc_hd__nor2_1
X_6141_ _6141_/A vssd1 vssd1 vccd1 vccd1 _6333_/D sky130_fd_sc_hd__clkbuf_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _4877_/B vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3284_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__inv_2
X_6072_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6308_/D sky130_fd_sc_hd__clkbuf_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5023_ _5023_/A _5023_/B vssd1 vssd1 vccd1 vccd1 _5024_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_674 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5925_ _6282_/Q _6293_/Q vssd1 vssd1 vccd1 vccd1 _5925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5856_ _5896_/S vssd1 vssd1 vccd1 vccd1 _5868_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4807_ _4798_/A _4798_/B _4801_/A vssd1 vssd1 vccd1 vccd1 _4812_/A sky130_fd_sc_hd__a21oi_4
X_5787_ _6241_/B _5787_/B vssd1 vssd1 vccd1 vccd1 _5787_/Y sky130_fd_sc_hd__nor2_1
X_4738_ _4738_/A _4738_/B _4738_/C vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__nor3_1
X_4669_ _4787_/B vssd1 vssd1 vccd1 vccd1 _4864_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6339_ _6359_/CLK _6339_/D vssd1 vssd1 vccd1 vccd1 _6339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6315__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_527 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5233__A2 _5355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_70 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6046__A _6061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3971_ _5158_/A _4210_/B vssd1 vssd1 vccd1 vccd1 _3972_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5710_ _5710_/A _5710_/B vssd1 vssd1 vccd1 vccd1 _5710_/X sky130_fd_sc_hd__xor2_2
XANTENNA__5885__A _5885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _5648_/A _5641_/B vssd1 vssd1 vccd1 vccd1 _5642_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5572_ _5572_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _5675_/B sky130_fd_sc_hd__xor2_4
XANTENNA__5932__B1 _5861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4523_ _4523_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__xor2_4
XANTENNA__5109__B _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3852__B _4088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4948__B _4961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4454_ _4565_/A _4565_/B vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__or2_1
X_4385_ _5325_/C vssd1 vssd1 vccd1 vccd1 _5511_/B sky130_fd_sc_hd__clkbuf_2
X_3405_ _6304_/Q vssd1 vssd1 vccd1 vccd1 _3405_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3336_ _3763_/A vssd1 vssd1 vccd1 vccd1 _4694_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6124_ _6124_/A vssd1 vssd1 vccd1 vccd1 _6327_/D sky130_fd_sc_hd__clkbuf_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A _6060_/C _6055_/C vssd1 vssd1 vccd1 vccd1 _6055_/X sky130_fd_sc_hd__and3_1
X_3267_ _3270_/A vssd1 vssd1 vccd1 vccd1 _3267_/Y sky130_fd_sc_hd__inv_2
X_5006_ _5006_/A _5006_/B vssd1 vssd1 vccd1 vccd1 _5016_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3198_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5908_ _5901_/A _5906_/B _5907_/X vssd1 vssd1 vccd1 vccd1 _5909_/B sky130_fd_sc_hd__o21a_1
X_5839_ _6378_/Q vssd1 vssd1 vccd1 vccd1 _5839_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5206__A2 _5489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_614 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__B1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4170_ _5404_/A _4207_/B _4167_/Y _4168_/X vssd1 vssd1 vccd1 vccd1 _4170_/X sky130_fd_sc_hd__a211o_1
XFILLER_96_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5174__D_N _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5850__C1 _6259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3954_ _5098_/A _4128_/B _4131_/B _5097_/A vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3885_ _4925_/A _4166_/B _3885_/C vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__and3_1
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5624_ _5624_/A _5624_/B vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__and2_1
X_5555_ _5585_/A _5585_/B _5554_/X vssd1 vssd1 vccd1 vccd1 _5562_/B sky130_fd_sc_hd__a21o_2
X_4506_ _4506_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4621_/B sky130_fd_sc_hd__xor2_4
X_5486_ _6275_/Q _5486_/B vssd1 vssd1 vccd1 vccd1 _5505_/C sky130_fd_sc_hd__and2_1
XFILLER_2_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4437_ _4438_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4558_/B sky130_fd_sc_hd__or2_1
XFILLER_116_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4368_ _4366_/A _4366_/B _4367_/X vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__a21oi_1
XFILLER_58_213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A io_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6107_ _6321_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6108_/A sky130_fd_sc_hd__and2_1
X_4299_ _5382_/A _4365_/B _4365_/C vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__and3_1
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3319_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_100_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6038_ _6036_/X _6042_/B _6023_/A vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__a21bo_1
XFILLER_66_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6563__79 vssd1 vssd1 vccd1 vccd1 _6563__79/HI _6563_/A sky130_fd_sc_hd__conb_1
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4883__B1 _4882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3670_ _3513_/A _3513_/B _3512_/A vssd1 vssd1 vccd1 vccd1 _3672_/C sky130_fd_sc_hd__a21o_1
XANTENNA__3683__A _5091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5363__A1 _5450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5340_ _5343_/B _5343_/A vssd1 vssd1 vccd1 vccd1 _5345_/A sky130_fd_sc_hd__and2b_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5271_ _5274_/A _5444_/B _5444_/C vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__and3_1
X_4222_ _4222_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4472_/B sky130_fd_sc_hd__and2_2
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4153_ _5294_/A _4153_/B _4153_/C vssd1 vssd1 vccd1 vccd1 _4188_/A sky130_fd_sc_hd__and3_1
X_4084_ _4126_/A _4126_/B _4083_/X vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__a21oi_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4961__B _4961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4986_ _4986_/A _4986_/B vssd1 vssd1 vccd1 vccd1 _4988_/C sky130_fd_sc_hd__xor2_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3937_ _4492_/A _3937_/B vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__and2_1
XFILLER_51_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3577__B _4882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3868_ _4051_/B vssd1 vssd1 vccd1 vccd1 _3906_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6587_ _6587_/A _3305_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_3799_ _5255_/A vssd1 vssd1 vccd1 vccd1 _5199_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5607_ _5675_/B _5608_/B vssd1 vssd1 vccd1 vccd1 _5613_/B sky130_fd_sc_hd__xnor2_1
X_5538_ _5590_/A _5590_/B _5537_/X vssd1 vssd1 vccd1 vccd1 _5586_/B sky130_fd_sc_hd__a21o_1
XFILLER_11_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5469_ _6275_/Q _5469_/B _5469_/C vssd1 vssd1 vccd1 vccd1 _5476_/B sky130_fd_sc_hd__and3_1
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5207__B _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6058__C1 _5904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _4840_/A _4840_/B _4840_/C vssd1 vssd1 vccd1 vccd1 _4852_/B sky130_fd_sc_hd__nand3_1
XANTENNA__3678__A _6280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6054__A _6060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4771_/A _4786_/A vssd1 vssd1 vccd1 vccd1 _4773_/B sky130_fd_sc_hd__nand2_1
X_6510_ _6510_/A _3216_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6527__46 vssd1 vssd1 vccd1 vccd1 _6527__46/HI _6527_/A sky130_fd_sc_hd__conb_1
X_3722_ _5007_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__and2_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3653_ _4815_/A _3653_/B _3653_/C vssd1 vssd1 vccd1 vccd1 _3693_/A sky130_fd_sc_hd__and3_2
X_6372_ _6375_/CLK _6372_/D vssd1 vssd1 vccd1 vccd1 _6372_/Q sky130_fd_sc_hd__dfxtp_1
X_5323_ _5323_/A _5323_/B vssd1 vssd1 vccd1 vccd1 _5333_/B sky130_fd_sc_hd__xor2_1
X_3584_ _3583_/A _3583_/C _3583_/B vssd1 vssd1 vccd1 vccd1 _3585_/C sky130_fd_sc_hd__a21oi_1
XFILLER_114_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5254_ _5257_/A _5257_/B vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__and2b_1
XFILLER_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4205_ _4237_/A _4204_/Y _4203_/A vssd1 vssd1 vccd1 vccd1 _4206_/B sky130_fd_sc_hd__a21oi_4
X_5185_ _5179_/A _5179_/B _5179_/C vssd1 vssd1 vccd1 vccd1 _5186_/D sky130_fd_sc_hd__a21o_1
X_4136_ _4139_/B _4139_/A vssd1 vssd1 vccd1 vccd1 _4141_/B sky130_fd_sc_hd__or2b_1
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4067_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4067_/X sky130_fd_sc_hd__and2b_1
XFILLER_83_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3822__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ _5109_/B vssd1 vssd1 vccd1 vccd1 _5145_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4882__A _4882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3945__B _4235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5941_ _5941_/A vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3201__A _3201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5872_ _6187_/A vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__clkbuf_2
X_4823_ _4823_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4835_/A sky130_fd_sc_hd__xor2_2
X_4754_ _4726_/B _4731_/B _3484_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _4755_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _3731_/A _3704_/C _3704_/A vssd1 vssd1 vccd1 vccd1 _3706_/C sky130_fd_sc_hd__a21o_1
X_4685_ _4687_/A _4687_/B vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__nand2_1
X_3636_ _4072_/A _4072_/B _4072_/C vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__a21o_1
X_6355_ _6357_/CLK _6355_/D vssd1 vssd1 vccd1 vccd1 _6355_/Q sky130_fd_sc_hd__dfxtp_1
X_3567_ _3566_/B _3567_/B vssd1 vssd1 vccd1 vccd1 _3567_/X sky130_fd_sc_hd__and2b_1
X_5306_ _5309_/B _5309_/A vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3871__A _4088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6286_ _6335_/CLK _6286_/D vssd1 vssd1 vccd1 vccd1 _6286_/Q sky130_fd_sc_hd__dfxtp_1
X_5237_ _5281_/A _5281_/B vssd1 vssd1 vccd1 vccd1 _5237_/Y sky130_fd_sc_hd__nor2_1
X_3498_ _3642_/A _3497_/B _3497_/C vssd1 vssd1 vccd1 vccd1 _3499_/C sky130_fd_sc_hd__a21o_1
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5168_ _5130_/A _5243_/B _5246_/B _5166_/A vssd1 vssd1 vccd1 vccd1 _5169_/B sky130_fd_sc_hd__a22oi_1
XFILLER_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4119_ _4119_/A _4167_/A _3940_/B vssd1 vssd1 vccd1 vccd1 _4122_/C sky130_fd_sc_hd__or3b_1
X_5099_ _5099_/A vssd1 vssd1 vccd1 vccd1 _5236_/B sky130_fd_sc_hd__clkbuf_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4207__A _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_274 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5181__C1 _4961_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5980__B _5980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__A1 _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _4518_/A _4518_/B _4469_/Y vssd1 vssd1 vccd1 vccd1 _4512_/B sky130_fd_sc_hd__a21bo_2
XFILLER_7_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3421_ _3645_/D vssd1 vssd1 vccd1 vccd1 _3692_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3352_ _4707_/A vssd1 vssd1 vccd1 vccd1 _4877_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6140_ _6140_/A input2/X vssd1 vssd1 vccd1 vccd1 _6141_/A sky130_fd_sc_hd__and2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__buf_6
XFILLER_97_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6071_ _6307_/Q _6073_/B vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__and2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5052_/A _5052_/B vssd1 vssd1 vccd1 vccd1 _5557_/A sky130_fd_sc_hd__nor2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _6282_/Q _6293_/Q vssd1 vssd1 vccd1 vccd1 _5924_/X sky130_fd_sc_hd__and2_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5855_ _5851_/X _5852_/Y _5853_/X _5854_/X vssd1 vssd1 vccd1 vccd1 _5896_/S sky130_fd_sc_hd__o22a_1
X_4806_ _4808_/B _4808_/A vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__or2b_1
X_5786_ _5838_/B _5786_/B vssd1 vssd1 vccd1 vccd1 _5787_/B sky130_fd_sc_hd__or2_1
X_4737_ _4738_/B _4738_/C _4738_/A vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__o21a_1
X_4668_ _3387_/A _5685_/A _6000_/A vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__a21o_1
X_3619_ _3619_/A _3619_/B vssd1 vssd1 vccd1 vccd1 _3619_/Y sky130_fd_sc_hd__nor2_1
X_6511__30 vssd1 vssd1 vccd1 vccd1 _6511__30/HI _6511_/A sky130_fd_sc_hd__conb_1
X_4599_ _4564_/Y _4571_/Y _4572_/Y _4578_/Y _4598_/X vssd1 vssd1 vccd1 vccd1 _4599_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6338_ _6359_/CLK _6338_/D vssd1 vssd1 vccd1 vccd1 _6338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6269_ _6382_/Q _6381_/Q _6269_/C vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__and3_1
XFILLER_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _4122_/B vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6569__85 vssd1 vssd1 vccd1 vccd1 _6569__85/HI _6569_/A sky130_fd_sc_hd__conb_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5640_ _5646_/A vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__clkbuf_2
X_5571_ _5571_/A _5571_/B vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4522_ _4522_/A _4522_/B vssd1 vssd1 vccd1 vccd1 _4624_/A sky130_fd_sc_hd__xnor2_2
X_4453_ _4451_/A _4451_/B _4575_/A vssd1 vssd1 vccd1 vccd1 _4565_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3404_ _6286_/Q _3549_/B _3549_/C vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__and3_1
X_4384_ _4384_/A _4384_/B vssd1 vssd1 vccd1 vccd1 _4459_/A sky130_fd_sc_hd__xnor2_1
X_3335_ _4664_/A vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6123_ _6326_/Q _6127_/B vssd1 vssd1 vccd1 vccd1 _6124_/A sky130_fd_sc_hd__and2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3266_ _3270_/A vssd1 vssd1 vccd1 vccd1 _3266_/Y sky130_fd_sc_hd__inv_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6060_/A _6060_/B vssd1 vssd1 vccd1 vccd1 _6055_/C sky130_fd_sc_hd__xnor2_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5005_ _4978_/A _4961_/B _4948_/C vssd1 vssd1 vccd1 vccd1 _5006_/B sky130_fd_sc_hd__a21oi_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _3201_/A vssd1 vssd1 vccd1 vccd1 _3197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6237__A _6259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5907_ _5755_/A _5899_/B _5902_/A vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _6379_/Q _5838_/B _5837_/Y vssd1 vssd1 vccd1 vccd1 _5838_/X sky130_fd_sc_hd__or3b_1
X_5769_ _6063_/A _6061_/A _5770_/A vssd1 vssd1 vccd1 vccd1 _5769_/X sky130_fd_sc_hd__and3b_1
XFILLER_108_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4414__A1 _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5914__A1 _3333_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_494 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _3840_/A _3785_/B _5885_/A vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _3875_/A _3875_/B _3883_/X vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__4305__A _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4169__B1 _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5905__A1 _5901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5623_ _5624_/A _5624_/B vssd1 vssd1 vccd1 vccd1 _5627_/B sky130_fd_sc_hd__xor2_1
X_5554_ _5554_/A _5554_/B _5554_/C vssd1 vssd1 vccd1 vccd1 _5554_/X sky130_fd_sc_hd__and3_1
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4505_ _4516_/A _4516_/B vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__nor2_1
X_5485_ _5485_/A _5485_/B _5504_/A vssd1 vssd1 vccd1 vccd1 _5488_/A sky130_fd_sc_hd__and3_1
XFILLER_105_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4436_ _4411_/A _4429_/Y _4433_/Y _4440_/B vssd1 vssd1 vccd1 vccd1 _4438_/B sky130_fd_sc_hd__o22a_1
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4367_ _5358_/A _4367_/B _4377_/B vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__and3_1
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _6106_/A vssd1 vssd1 vccd1 vccd1 _6321_/D sky130_fd_sc_hd__clkbuf_1
X_3318_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3318_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4298_ _6276_/Q vssd1 vssd1 vccd1 vccd1 _5382_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3249_/Y sky130_fd_sc_hd__inv_2
X_6037_ _6036_/B _6036_/C _6036_/A vssd1 vssd1 vccd1 vccd1 _6042_/B sky130_fd_sc_hd__o21ai_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539__55 vssd1 vssd1 vccd1 vccd1 _6539__55/HI _6539_/A sky130_fd_sc_hd__conb_1
XANTENNA__5363__A2 _5485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5270_ _5270_/A vssd1 vssd1 vccd1 vccd1 _5444_/C sky130_fd_sc_hd__clkbuf_2
X_4221_ _4224_/A _4224_/B vssd1 vssd1 vccd1 vccd1 _4222_/B sky130_fd_sc_hd__or2b_1
XFILLER_102_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _5165_/A _4412_/B _4153_/C _5208_/A vssd1 vssd1 vccd1 vccd1 _4188_/B sky130_fd_sc_hd__a22oi_2
XFILLER_110_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4083_ _4078_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__and2b_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3204__A _3208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4985_ _5619_/A _4994_/B vssd1 vssd1 vccd1 vccd1 _4986_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3936_ _4482_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _3937_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3867_ _3883_/A _3867_/B vssd1 vssd1 vccd1 vccd1 _3875_/A sky130_fd_sc_hd__xnor2_1
X_3798_ _5320_/A vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__clkbuf_2
X_6586_ _6586_/A _3304_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_5606_ _5606_/A _5606_/B vssd1 vssd1 vccd1 vccd1 _5608_/B sky130_fd_sc_hd__xnor2_1
X_5537_ _5408_/B _5537_/B vssd1 vssd1 vccd1 vccd1 _5537_/X sky130_fd_sc_hd__and2b_1
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6587__103 vssd1 vssd1 vccd1 vccd1 _6587__103/HI _6587_/A sky130_fd_sc_hd__conb_1
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5468_ _5468_/A _5493_/A vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__nor2_1
X_4419_ _4426_/A _4426_/B vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__and2_1
X_5399_ _5421_/A _5421_/B _5397_/A vssd1 vssd1 vccd1 vccd1 _5401_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5207__C _5469_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6230__B1 _5952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4770_ _4771_/A _4770_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _4786_/A sky130_fd_sc_hd__nand3_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3721_ _4122_/B vssd1 vssd1 vccd1 vccd1 _4235_/B sky130_fd_sc_hd__clkbuf_2
X_3652_ _3690_/A _3652_/B _3652_/C vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__and3_1
X_6371_ _6375_/CLK _6371_/D vssd1 vssd1 vccd1 vccd1 _6371_/Q sky130_fd_sc_hd__dfxtp_1
X_3583_ _3583_/A _3583_/B _3583_/C vssd1 vssd1 vccd1 vccd1 _3585_/B sky130_fd_sc_hd__and3_1
X_5322_ _5322_/A _5322_/B vssd1 vssd1 vccd1 vccd1 _5323_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5253_ _5286_/A _5286_/B _5252_/A vssd1 vssd1 vccd1 vccd1 _5257_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4204_ _4237_/B vssd1 vssd1 vccd1 vccd1 _4204_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5184_ _4059_/A _5183_/B _5183_/C _5183_/D vssd1 vssd1 vccd1 vccd1 _5186_/C sky130_fd_sc_hd__a22o_1
X_4135_ _4143_/A _4143_/B _4134_/X vssd1 vssd1 vccd1 vccd1 _4139_/A sky130_fd_sc_hd__a21o_1
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5133__B _5172_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4066_/A _4066_/B vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4968_ _4954_/Y _4966_/X _4967_/Y _4951_/Y vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _3919_/A _3919_/B _3919_/C vssd1 vssd1 vccd1 vccd1 _3920_/B sky130_fd_sc_hd__and3_1
X_4899_ _4726_/A _3632_/C _4905_/A _4898_/Y vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__o22ai_2
XANTENNA__5308__B _5308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6569_ _6569_/A _3285_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_105_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3510__A1 _3536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5978__B _5980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5234__A _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6065__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _5940_/A _5941_/A vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__xnor2_1
XFILLER_92_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5871_ _6098_/A vssd1 vssd1 vccd1 vccd1 _6187_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4822_ _4822_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4838_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4753_ _4664_/A _4764_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__a21o_1
X_3704_ _3704_/A _3731_/A _3704_/C vssd1 vssd1 vccd1 vccd1 _3731_/B sky130_fd_sc_hd__nand3_1
X_4684_ _4736_/A _4736_/B _4683_/A vssd1 vssd1 vccd1 vccd1 _4687_/B sky130_fd_sc_hd__o21ai_1
X_3635_ _4110_/B _3635_/B vssd1 vssd1 vccd1 vccd1 _4072_/C sky130_fd_sc_hd__nand2_1
X_6354_ _6357_/CLK _6354_/D vssd1 vssd1 vccd1 vccd1 _6354_/Q sky130_fd_sc_hd__dfxtp_1
X_3566_ _3567_/B _3566_/B vssd1 vssd1 vccd1 vccd1 _3570_/B sky130_fd_sc_hd__xnor2_1
X_5305_ _5309_/A _5309_/B vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__and2b_1
X_3497_ _3642_/A _3497_/B _3497_/C vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__nand3_1
X_6285_ _6359_/CLK _6285_/D vssd1 vssd1 vccd1 vccd1 _6285_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5236_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _5281_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5167_ _5382_/B _5382_/C vssd1 vssd1 vccd1 vccd1 _5246_/B sky130_fd_sc_hd__and2_1
XFILLER_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4118_ _5231_/B _4268_/B vssd1 vssd1 vccd1 vccd1 _4167_/A sky130_fd_sc_hd__nand2_2
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5098_ _5098_/A _5099_/A _5098_/C vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__and3_1
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4049_ _5355_/A vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_359 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5038__B _5038_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5181__B1 _4062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3302__A _3306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_60 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3420_ _3458_/A _4707_/B vssd1 vssd1 vccd1 vccd1 _3645_/D sky130_fd_sc_hd__xor2_1
XANTENNA__4787__B _4787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3351_ _3522_/A vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3282_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__inv_2
X_6070_ _6070_/A vssd1 vssd1 vccd1 vccd1 _6307_/D sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5021_ _5050_/A _5050_/B _5020_/A vssd1 vssd1 vccd1 vccd1 _5052_/B sky130_fd_sc_hd__o21a_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3212__A _3214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5923_ _5936_/A vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5854_ _6314_/Q _6323_/Q vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__and2b_1
X_4805_ _4805_/A _4805_/B vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__xor2_2
X_5785_ _5719_/Y _5690_/A _5815_/B _5717_/Y _5784_/Y vssd1 vssd1 vccd1 vccd1 _5786_/B
+ sky130_fd_sc_hd__o221a_1
X_4736_ _4736_/A _4736_/B vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__xor2_1
XFILLER_107_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4667_ _4644_/A _4664_/X _4666_/X vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__a21boi_1
XFILLER_107_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3618_ _3627_/B _3627_/C _3627_/A vssd1 vssd1 vccd1 vccd1 _3626_/B sky130_fd_sc_hd__a21bo_1
X_4598_ _4572_/Y _4578_/Y _4584_/Y _4585_/Y _4597_/X vssd1 vssd1 vccd1 vccd1 _4598_/X
+ sky130_fd_sc_hd__a221o_1
X_6337_ _6345_/CLK _6337_/D vssd1 vssd1 vccd1 vccd1 _6337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3549_ _6285_/Q _3549_/B _3549_/C vssd1 vssd1 vccd1 vccd1 _3575_/C sky130_fd_sc_hd__and3_1
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4269__A2 _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6268_ _6381_/Q _6269_/C _6267_/Y vssd1 vssd1 vccd1 vccd1 _6381_/D sky130_fd_sc_hd__o21a_1
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _4059_/A _5218_/D _5216_/X _5217_/Y vssd1 vssd1 vccd1 vccd1 _5221_/C sky130_fd_sc_hd__o2bb2a_1
X_6199_ _6356_/Q _6201_/B vssd1 vssd1 vccd1 vccd1 _6200_/A sky130_fd_sc_hd__and2_1
XANTENNA__5602__A _5737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_112 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5570_ _5579_/A _5570_/B vssd1 vssd1 vccd1 vccd1 _5572_/A sky130_fd_sc_hd__and2_1
X_4521_ _4521_/A _4521_/B vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__or2_1
XFILLER_116_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4452_ _4574_/A _4574_/B vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3403_ _3400_/X _4749_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _3549_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__3207__A _3208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4383_ _4461_/B _4383_/B vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__xnor2_2
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6122_ _6122_/A vssd1 vssd1 vccd1 vccd1 _6326_/D sky130_fd_sc_hd__clkbuf_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _6290_/Q vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3265_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3270_/A sky130_fd_sc_hd__buf_6
XFILLER_105_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6061_/B _6023_/X _6052_/X _5904_/X vssd1 vssd1 vccd1 vccd1 _6302_/D sky130_fd_sc_hd__o211a_1
X_5004_ _5004_/A _5004_/B vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__xor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3196_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3201_/A sky130_fd_sc_hd__buf_6
XFILLER_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6384__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5906_ _5906_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__xor2_1
XFILLER_22_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5837_ _5717_/Y _5690_/B _5773_/B _5719_/Y _5836_/Y vssd1 vssd1 vccd1 vccd1 _5837_/Y
+ sky130_fd_sc_hd__o221ai_2
X_5768_ _6367_/Q _5697_/Y _5708_/X _5764_/X _6259_/A vssd1 vssd1 vccd1 vccd1 _6538_/A
+ sky130_fd_sc_hd__a221oi_4
X_4719_ _4719_/A _4719_/B _4719_/C vssd1 vssd1 vccd1 vccd1 _4720_/B sky130_fd_sc_hd__nand3_1
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5699_ _5819_/A _5699_/B vssd1 vssd1 vccd1 vccd1 _5741_/B sky130_fd_sc_hd__or2_1
XFILLER_107_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5687__A1 _6061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4414__A2 _4153_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6163__A _6187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_50 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3952_ _4386_/A vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__buf_4
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ _3883_/A _3867_/B vssd1 vssd1 vccd1 vccd1 _3883_/X sky130_fd_sc_hd__or2b_1
XANTENNA__4305__B _4337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5622_ _5622_/A _5622_/B vssd1 vssd1 vccd1 vccd1 _5624_/B sky130_fd_sc_hd__and2_1
X_5553_ _5589_/A _5589_/B _5552_/X vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__a21o_1
X_4504_ _4546_/A _4546_/B vssd1 vssd1 vccd1 vccd1 _4516_/B sky130_fd_sc_hd__nand2_1
X_5484_ _5484_/A _5484_/B _5484_/C vssd1 vssd1 vccd1 vccd1 _5504_/A sky130_fd_sc_hd__and3_1
X_4435_ _4435_/A _4435_/B vssd1 vssd1 vccd1 vccd1 _4440_/B sky130_fd_sc_hd__or2_1
X_4366_ _4366_/A _4366_/B vssd1 vssd1 vccd1 vccd1 _4377_/B sky130_fd_sc_hd__xor2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3317_/Y sky130_fd_sc_hd__inv_2
X_6105_ _6320_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6106_/A sky130_fd_sc_hd__and2_1
X_4297_ _4297_/A _4297_/B vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__xnor2_2
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3248_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3248_/Y sky130_fd_sc_hd__inv_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6036_/A _6036_/B _6036_/C vssd1 vssd1 vccd1 vccd1 _6036_/X sky130_fd_sc_hd__or3_1
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4109__C _4365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3310__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5348__B1 _5489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4571__A1 _4569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4220_ _4220_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4224_/B sky130_fd_sc_hd__xnor2_2
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4151_ _4410_/B vssd1 vssd1 vccd1 vccd1 _4153_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4082_ _4082_/A _4082_/B vssd1 vssd1 vccd1 vccd1 _4126_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _4998_/A _4998_/B _4998_/C vssd1 vssd1 vccd1 vccd1 _5023_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3220__A _3220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ _4496_/A _3935_/B vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__and2_1
X_3866_ _3892_/B _3866_/B vssd1 vssd1 vccd1 vccd1 _3867_/B sky130_fd_sc_hd__nor2_1
X_5605_ _5605_/A vssd1 vssd1 vccd1 vccd1 _5605_/Y sky130_fd_sc_hd__inv_2
X_3797_ _4266_/A vssd1 vssd1 vccd1 vccd1 _5320_/A sky130_fd_sc_hd__clkbuf_2
X_6585_ _6585_/A _3303_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XANTENNA__4051__A _4059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4562__A1 _5627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5536_ _5598_/A _5598_/B _5535_/Y vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__a21bo_1
XFILLER_105_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5467_ _5468_/A _6276_/Q _5505_/B _5491_/A vssd1 vssd1 vccd1 vccd1 _5493_/A sky130_fd_sc_hd__and4b_1
X_4418_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4426_/B sky130_fd_sc_hd__xnor2_1
X_5398_ _5398_/A _5398_/B vssd1 vssd1 vccd1 vccd1 _5421_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4349_ _4369_/A _4369_/B _4348_/Y vssd1 vssd1 vccd1 vccd1 _4354_/B sky130_fd_sc_hd__o21a_1
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6019_ _6020_/A _6020_/B vssd1 vssd1 vccd1 vccd1 _6019_/X sky130_fd_sc_hd__or2_1
XFILLER_100_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6058__A1 _6061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3305__A _3306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_84 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3720_ _3782_/A _3720_/B vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _3661_/A _3733_/A vssd1 vssd1 vccd1 vccd1 _3688_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6370_ _6375_/CLK _6370_/D vssd1 vssd1 vccd1 vccd1 _6370_/Q sky130_fd_sc_hd__dfxtp_1
X_3582_ _3564_/A _3563_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3583_/C sky130_fd_sc_hd__a21o_1
X_5321_ _5321_/A _5321_/B vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3499__A_N _3476_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5252_ _5252_/A _5252_/B vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4203_ _4203_/A _4203_/B vssd1 vssd1 vccd1 vccd1 _4237_/B sky130_fd_sc_hd__or2_1
X_5183_ _5183_/A _5183_/B _5183_/C _5183_/D vssd1 vssd1 vccd1 vccd1 _5186_/B sky130_fd_sc_hd__nand4_2
X_4134_ _4127_/B _4134_/B vssd1 vssd1 vccd1 vccd1 _4134_/X sky130_fd_sc_hd__and2b_1
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4065_ _4009_/B _4057_/X _4056_/Y _4041_/X vssd1 vssd1 vccd1 vccd1 _4066_/B sky130_fd_sc_hd__a211oi_1
XFILLER_71_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4967_ _4694_/B _4933_/B _4950_/Y _4953_/A vssd1 vssd1 vccd1 vccd1 _4967_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3918_ _3919_/A _3919_/B _3919_/C vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__a21oi_1
X_4898_ _4898_/A _4898_/B vssd1 vssd1 vccd1 vccd1 _4898_/Y sky130_fd_sc_hd__nor2_1
X_6518__37 vssd1 vssd1 vccd1 vccd1 _6518__37/HI _6518_/A sky130_fd_sc_hd__conb_1
X_3849_ _5134_/A vssd1 vssd1 vccd1 vccd1 _5098_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_674 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6568_ _6568_/A _3284_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_98_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5519_ _5519_/A _5519_/B vssd1 vssd1 vccd1 vccd1 _5520_/A sky130_fd_sc_hd__or2_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6499_ _6499_/A _3201_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5605__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6532__51 vssd1 vssd1 vccd1 vccd1 _6532__51/HI _6532_/A sky130_fd_sc_hd__conb_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__B _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5870_ _5980_/B vssd1 vssd1 vccd1 vccd1 _6098_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4821_ _4830_/B _4856_/A vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__and2b_1
XFILLER_61_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _3690_/A _4751_/X _4757_/A vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__a21bo_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4683_ _4683_/A _4683_/B vssd1 vssd1 vccd1 vccd1 _4736_/B sky130_fd_sc_hd__nand2_1
X_3703_ _3739_/B _3702_/C _3702_/A vssd1 vssd1 vccd1 vccd1 _3704_/C sky130_fd_sc_hd__a21o_1
X_3634_ _3633_/X _3634_/B vssd1 vssd1 vccd1 vccd1 _3635_/B sky130_fd_sc_hd__and2b_1
X_6353_ _6357_/CLK _6353_/D vssd1 vssd1 vccd1 vccd1 _6353_/Q sky130_fd_sc_hd__dfxtp_1
X_3565_ _3565_/A _3565_/B vssd1 vssd1 vccd1 vccd1 _3566_/B sky130_fd_sc_hd__xnor2_1
X_5304_ _5259_/B _5283_/X _5302_/B _5303_/Y vssd1 vssd1 vccd1 vccd1 _5309_/B sky130_fd_sc_hd__o31a_1
X_3496_ _3496_/A _3661_/C vssd1 vssd1 vccd1 vccd1 _3497_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6284_ _6359_/CLK _6284_/D vssd1 vssd1 vccd1 vccd1 _6284_/Q sky130_fd_sc_hd__dfxtp_1
X_5235_ _5235_/A _5235_/B vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5166_ _5166_/A _5274_/D _5166_/C vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__and3_1
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4117_ _4117_/A _4117_/B vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__xnor2_1
X_5097_ _5097_/A _5134_/B vssd1 vssd1 vccd1 vccd1 _5098_/C sky130_fd_sc_hd__and2_1
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4048_ _5278_/A vssd1 vssd1 vccd1 vccd1 _5355_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5999_ _6000_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6001_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4504__A _4546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5953__B1 _5952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6290__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_302 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ _6286_/Q vssd1 vssd1 vccd1 vccd1 _3522_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5020_ _5020_/A _5020_/B vssd1 vssd1 vccd1 vccd1 _5050_/B sky130_fd_sc_hd__nand2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3281_/Y sky130_fd_sc_hd__inv_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__B2 _6291_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5922_ _5922_/A vssd1 vssd1 vccd1 vccd1 _6283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5853_ _6323_/Q _6314_/Q vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__and2b_1
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4324__A _5355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4804_ _4802_/A _4802_/B _4803_/X vssd1 vssd1 vccd1 vccd1 _4808_/B sky130_fd_sc_hd__o21a_1
XFILLER_61_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5784_ _5715_/A _5777_/B _5841_/B vssd1 vssd1 vccd1 vccd1 _5784_/Y sky130_fd_sc_hd__a21oi_1
X_4735_ _4761_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4738_/C sky130_fd_sc_hd__nor2_1
XFILLER_9_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4666_ _4664_/A _4864_/D _4785_/C _4820_/A vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__a22o_1
X_4597_ _4589_/X _4596_/X _4584_/Y _4585_/Y vssd1 vssd1 vccd1 vccd1 _4597_/X sky130_fd_sc_hd__o2bb2a_1
X_3617_ _3617_/A _3617_/B _3617_/C vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__nand3_1
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6336_ _6345_/CLK _6336_/D vssd1 vssd1 vccd1 vccd1 _6336_/Q sky130_fd_sc_hd__dfxtp_1
X_3548_ _3548_/A _3576_/A vssd1 vssd1 vccd1 vccd1 _3552_/A sky130_fd_sc_hd__and2_1
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4994__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3479_ _3479_/A vssd1 vssd1 vccd1 vccd1 _3645_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5466__A2 _4370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6267_ _6267_/A _6267_/B vssd1 vssd1 vccd1 vccd1 _6267_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5218_ _5216_/X _5217_/Y _5236_/A _5218_/D vssd1 vssd1 vccd1 vccd1 _5221_/B sky130_fd_sc_hd__and4bb_1
XFILLER_57_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6198_ _6198_/A vssd1 vssd1 vccd1 vccd1 _6356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5149_ _5113_/A _5113_/C _5113_/B vssd1 vssd1 vccd1 vccd1 _5149_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6502__21 vssd1 vssd1 vccd1 vccd1 _6502__21/HI _6502_/A sky130_fd_sc_hd__conb_1
XFILLER_109_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5231__C _5273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4520_ _4537_/A _4536_/A _4536_/B _4017_/A vssd1 vssd1 vccd1 vccd1 _4522_/A sky130_fd_sc_hd__a31o_1
XFILLER_116_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4451_ _4451_/A _4451_/B vssd1 vssd1 vccd1 vccd1 _4574_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3402_ _3386_/A _3391_/A _6298_/Q vssd1 vssd1 vccd1 vccd1 _4769_/B sky130_fd_sc_hd__a21o_2
X_4382_ _4384_/A _4384_/B _4381_/X vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__o21ba_1
X_6121_ _6325_/Q _6127_/B vssd1 vssd1 vccd1 vccd1 _6122_/A sky130_fd_sc_hd__and2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _5613_/A vssd1 vssd1 vccd1 vccd1 _3333_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3264_ input1/X vssd1 vssd1 vccd1 vccd1 _3289_/A sky130_fd_sc_hd__buf_2
XFILLER_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6050_/X _6060_/C _6023_/A vssd1 vssd1 vccd1 vccd1 _6052_/X sky130_fd_sc_hd__a21bo_1
X_5003_ _5003_/A _5003_/B vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__xnor2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3223__A _3226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3195_ _3195_/A vssd1 vssd1 vccd1 vccd1 _3195_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5905_ _5901_/A _5910_/A _5902_/X _5903_/Y _5904_/X vssd1 vssd1 vccd1 vccd1 _6279_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5836_ _5715_/A _5819_/B _5777_/A vssd1 vssd1 vccd1 vccd1 _5836_/Y sky130_fd_sc_hd__a21oi_1
X_5767_ _6270_/A vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__clkbuf_4
X_4718_ _4718_/A _4718_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__xor2_1
X_5698_ _5698_/A vssd1 vssd1 vccd1 vccd1 _5906_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4649_ _4656_/B _4645_/Y _4648_/X vssd1 vssd1 vccd1 vccd1 _4680_/B sky130_fd_sc_hd__o21ba_1
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6319_ _6369_/CLK _6319_/D vssd1 vssd1 vccd1 vccd1 _6319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6163__B input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3925__A2 _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6574__90 vssd1 vssd1 vccd1 vccd1 _6574__90/HI _6574_/A sky130_fd_sc_hd__conb_1
XANTENNA__3308__A _3312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _6277_/Q vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__inv_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3882_ _3965_/B _3965_/A vssd1 vssd1 vccd1 vccd1 _3938_/B sky130_fd_sc_hd__or2b_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4305__C _4337_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ _5621_/A _5621_/B _5629_/A vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__or3_1
XANTENNA__4602__A _4621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5552_ _5120_/B _5552_/B vssd1 vssd1 vccd1 vccd1 _5552_/X sky130_fd_sc_hd__and2b_1
X_4503_ _4509_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4546_/B sky130_fd_sc_hd__o21ai_2
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3218__A _3220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5483_ _5483_/A _5483_/B vssd1 vssd1 vccd1 vccd1 _5497_/A sky130_fd_sc_hd__xnor2_1
X_4434_ _5349_/A _4580_/B _5484_/B vssd1 vssd1 vccd1 vccd1 _4435_/B sky130_fd_sc_hd__a21oi_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ _5416_/A _4365_/B _4365_/C vssd1 vssd1 vccd1 vccd1 _4366_/B sky130_fd_sc_hd__and3_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _6104_/A vssd1 vssd1 vccd1 vccd1 _6320_/D sky130_fd_sc_hd__clkbuf_1
X_6493__12 vssd1 vssd1 vccd1 vccd1 _6493__12/HI _6493_/A sky130_fd_sc_hd__conb_1
X_3316_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3316_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4296_ _4296_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4465_/B sky130_fd_sc_hd__xnor2_4
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6026_/B _6035_/B vssd1 vssd1 vccd1 vccd1 _6036_/C sky130_fd_sc_hd__and2b_1
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4049__A _5355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3247_ _3251_/A vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__inv_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_606 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5819_ _5819_/A _5819_/B vssd1 vssd1 vccd1 vccd1 _5820_/A sky130_fd_sc_hd__or2_1
XFILLER_10_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5608__A _5675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5293__B1 _5505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4150_ _4301_/B vssd1 vssd1 vccd1 vccd1 _4410_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4081_ _4089_/A _4089_/B vssd1 vssd1 vccd1 vccd1 _4082_/B sky130_fd_sc_hd__xor2_1
XFILLER_68_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3501__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4983_ _4983_/A _4991_/B vssd1 vssd1 vccd1 vccd1 _4998_/C sky130_fd_sc_hd__xnor2_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3934_ _3934_/A _3934_/B vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3865_ _4960_/A _4138_/B _3864_/C vssd1 vssd1 vccd1 vccd1 _3866_/B sky130_fd_sc_hd__a21oi_1
X_5604_ _5676_/A _5610_/B vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__xnor2_1
X_6584_ _6584_/A _3302_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_3796_ _5349_/A vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4051__B _4051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5535_ _5535_/A _5535_/B vssd1 vssd1 vccd1 vccd1 _5535_/Y sky130_fd_sc_hd__nand2_1
X_5466_ _5440_/A _4370_/B _5440_/C vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__a21o_1
X_4417_ _4417_/A _4417_/B vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__nor2_1
X_5397_ _5397_/A _5397_/B vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6259__A _6259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_A io_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4348_ _4348_/A _4348_/B vssd1 vssd1 vccd1 vccd1 _4348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4279_ _6281_/Q _4279_/B vssd1 vssd1 vccd1 vccd1 _4280_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _6006_/X _6011_/B _6009_/B vssd1 vssd1 vccd1 vccd1 _6020_/B sky130_fd_sc_hd__o21a_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_650 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6544__60 vssd1 vssd1 vccd1 vccd1 _6544__60/HI _6544_/A sky130_fd_sc_hd__conb_1
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3321__A _3321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3650_ _3649_/B _3649_/C _3649_/A vssd1 vssd1 vccd1 vccd1 _3657_/B sky130_fd_sc_hd__a21o_1
X_3581_ _3594_/A _3594_/B _3595_/B _3580_/Y vssd1 vssd1 vccd1 vccd1 _3583_/B sky130_fd_sc_hd__a31o_1
X_5320_ _5320_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5321_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _5251_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__or2_1
X_4202_ _4201_/B _4202_/B vssd1 vssd1 vccd1 vccd1 _4203_/B sky130_fd_sc_hd__and2b_1
X_5182_ _4053_/A _5218_/D _5174_/A _5180_/X vssd1 vssd1 vccd1 vccd1 _5183_/D sky130_fd_sc_hd__a211o_1
XFILLER_68_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4133_ _4133_/A _4138_/C vssd1 vssd1 vccd1 vccd1 _4143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _5866_/A _4484_/B _4055_/B _4063_/X vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__a31oi_4
XANTENNA__3231__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4232__A1 _4059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3885__B _4166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4966_ _4966_/A _4957_/B vssd1 vssd1 vccd1 vccd1 _4966_/X sky130_fd_sc_hd__or2b_1
X_3917_ _3934_/A _3917_/B vssd1 vssd1 vccd1 vccd1 _3919_/C sky130_fd_sc_hd__nand2_1
X_4897_ _4897_/A _4897_/B vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__or2_1
XFILLER_20_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4062__A _4062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3848_ _5195_/A vssd1 vssd1 vccd1 vccd1 _5134_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6567_ _6567_/A _3282_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_3779_ _3715_/A _3747_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5518_ _5514_/A _5514_/C _5514_/B vssd1 vssd1 vccd1 vccd1 _5521_/A sky130_fd_sc_hd__a21boi_1
X_6498_ _6498_/A _3200_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5449_ _5449_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3316__A _3318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4147__A _4340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4820_ _4820_/A _4820_/B vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__nand2_2
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4751_ _4815_/A _4879_/D _4787_/C vssd1 vssd1 vccd1 vccd1 _4751_/X sky130_fd_sc_hd__and3_1
XANTENNA__5962__A1 _5957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4682_ _4682_/A _4682_/B _4682_/C vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__nand3_1
X_3702_ _3702_/A _3739_/B _3702_/C vssd1 vssd1 vccd1 vccd1 _3731_/A sky130_fd_sc_hd__nand3_1
X_3633_ _3633_/A _3632_/X vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__or2b_1
XFILLER_108_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6352_ _6384_/CLK _6352_/D vssd1 vssd1 vccd1 vccd1 _6352_/Q sky130_fd_sc_hd__dfxtp_1
X_3564_ _3564_/A _3583_/A vssd1 vssd1 vccd1 vccd1 _3567_/B sky130_fd_sc_hd__nand2_1
X_5303_ _5339_/A _5339_/B vssd1 vssd1 vccd1 vccd1 _5303_/Y sky130_fd_sc_hd__nand2_1
X_3495_ _3495_/A _3495_/B vssd1 vssd1 vccd1 vccd1 _3661_/C sky130_fd_sc_hd__xnor2_1
X_6283_ _6384_/CLK _6283_/D vssd1 vssd1 vccd1 vccd1 _6283_/Q sky130_fd_sc_hd__dfxtp_1
X_5234_ _5404_/A _5278_/B vssd1 vssd1 vccd1 vccd1 _5235_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3226__A _3226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5165_ _5165_/A _5471_/B _5471_/C vssd1 vssd1 vccd1 vccd1 _5166_/C sky130_fd_sc_hd__and3_1
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ _4114_/A _4153_/B _4156_/A vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__a21oi_2
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5096_ _5070_/B _5091_/Y _5123_/A _5123_/B vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__o22ai_2
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4047_ _5358_/A vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _6000_/B vssd1 vssd1 vccd1 vccd1 _6016_/B sky130_fd_sc_hd__clkbuf_1
X_4949_ _4947_/A _4947_/B _5006_/A vssd1 vssd1 vccd1 vccd1 _4972_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__4504__B _4546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5953__A1 _5955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5616__A _5672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3280_ _3282_/A vssd1 vssd1 vccd1 vccd1 _3280_/Y sky130_fd_sc_hd__inv_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5921_ _6323_/Q _6073_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__and2_1
XFILLER_81_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_594 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ _6384_/Q _6283_/Q vssd1 vssd1 vccd1 vccd1 _5852_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6092__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4324__B _4324_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4803_ _4823_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__or2_1
XFILLER_21_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5783_ _6371_/Q vssd1 vssd1 vccd1 vccd1 _6241_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4734_ _4738_/B _4734_/B vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__or2_2
XFILLER_9_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4665_ _4769_/B vssd1 vssd1 vccd1 vccd1 _4785_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4596_ _5866_/A _4595_/B _4594_/X _4595_/Y _4589_/A vssd1 vssd1 vccd1 vccd1 _4596_/X
+ sky130_fd_sc_hd__a32o_1
X_3616_ _3629_/B _3614_/Y _3629_/A vssd1 vssd1 vccd1 vccd1 _3627_/C sky130_fd_sc_hd__o21a_1
X_6335_ _6335_/CLK _6335_/D vssd1 vssd1 vccd1 vccd1 _6335_/Q sky130_fd_sc_hd__dfxtp_1
X_3547_ _6286_/Q _3547_/B vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__and2_1
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6266_ _6381_/Q _6269_/C vssd1 vssd1 vccd1 vccd1 _6267_/B sky130_fd_sc_hd__and2_1
X_3478_ _4651_/A _3601_/B _3446_/D _3477_/X vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__a31o_1
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5217_ _4323_/A _5013_/B _5198_/A _5215_/X vssd1 vssd1 vccd1 vccd1 _5217_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6197_ _6355_/Q _6197_/B vssd1 vssd1 vccd1 vccd1 _6198_/A sky130_fd_sc_hd__and2_1
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5148_ _5141_/X _5151_/B _5148_/C _5148_/D vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__and4b_1
X_5079_ _5114_/B _5114_/C _5114_/A vssd1 vssd1 vccd1 vccd1 _5083_/B sky130_fd_sc_hd__a21boi_2
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5346__A _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5862__B1 _5861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4450_ _5865_/A _5511_/B _4587_/A _4581_/B vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__or4_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4381_ _4380_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4381_/X sky130_fd_sc_hd__and2b_1
X_3401_ _3401_/A vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6120_ _6120_/A vssd1 vssd1 vccd1 vccd1 _6325_/D sky130_fd_sc_hd__clkbuf_1
X_3332_ _5605_/A vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__clkbuf_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3263_/A vssd1 vssd1 vccd1 vccd1 _3263_/Y sky130_fd_sc_hd__inv_2
X_6051_ _6051_/A _6050_/A vssd1 vssd1 vccd1 vccd1 _6060_/C sky130_fd_sc_hd__or2b_1
X_5002_ _5004_/A _5004_/B vssd1 vssd1 vccd1 vccd1 _5050_/A sky130_fd_sc_hd__or2_1
X_3194_ _3195_/A vssd1 vssd1 vccd1 vccd1 _3194_/Y sky130_fd_sc_hd__inv_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5904_ _6201_/B vssd1 vssd1 vccd1 vccd1 _5904_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5908__A1 _5901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5835_ _6378_/Q _5827_/Y _5829_/X _5833_/X _5834_/X vssd1 vssd1 vccd1 vccd1 _5835_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5766_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4717_ _5966_/A _4814_/B vssd1 vssd1 vccd1 vccd1 _4718_/B sky130_fd_sc_hd__nor2_1
X_5697_ _3333_/X _3384_/X _5696_/X vssd1 vssd1 vccd1 vccd1 _5697_/Y sky130_fd_sc_hd__o21ai_2
X_4648_ _4656_/B _4647_/Y _4645_/Y vssd1 vssd1 vccd1 vccd1 _4648_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4579_ _5865_/A _5511_/B vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6318_ _6369_/CLK _6318_/D vssd1 vssd1 vccd1 vccd1 _6318_/Q sky130_fd_sc_hd__dfxtp_1
X_6249_ _6267_/A _6249_/B vssd1 vssd1 vccd1 vccd1 _6249_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3950_ _3950_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _3956_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ _3881_/A _3881_/B vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__xor2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_364 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5620_ _5627_/A vssd1 vssd1 vccd1 vccd1 _5755_/A sky130_fd_sc_hd__clkbuf_2
X_5551_ _5596_/B _5597_/B _5550_/X vssd1 vssd1 vccd1 vccd1 _5589_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4502_ _4509_/A _4502_/B _4502_/C vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__or3_2
X_5482_ _5482_/A _5482_/B vssd1 vssd1 vccd1 vccd1 _5500_/A sky130_fd_sc_hd__xnor2_1
X_4433_ _4440_/A vssd1 vssd1 vccd1 vccd1 _4433_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5714__A _5714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4364_ _6275_/Q vssd1 vssd1 vccd1 vccd1 _5416_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4295_ _4467_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__xor2_4
XFILLER_112_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6319_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6104_/A sky130_fd_sc_hd__and2_1
X_3315_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3315_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3246_ _3258_/A vssd1 vssd1 vccd1 vccd1 _3251_/A sky130_fd_sc_hd__buf_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6299_/Q _6016_/A _6060_/B vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__o21a_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6251__B1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5818_ _3333_/X _3384_/X _5817_/X vssd1 vssd1 vccd1 vccd1 _5818_/Y sky130_fd_sc_hd__o21ai_2
X_5749_ _5749_/A _5749_/B vssd1 vssd1 vccd1 vccd1 _5749_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5624__A _5624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5348__A2 _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3319__A _3321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4080_ _5133_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4089_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6233__B1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4982_ _4975_/A _4963_/B _4981_/X vssd1 vssd1 vccd1 vccd1 _4991_/B sky130_fd_sc_hd__o21ai_1
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3933_ _3934_/A _3934_/B vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__or2_2
X_3864_ _3903_/A _4138_/B _3864_/C vssd1 vssd1 vccd1 vccd1 _3892_/B sky130_fd_sc_hd__and3_1
X_5603_ _5603_/A _5603_/B vssd1 vssd1 vccd1 vccd1 _5610_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__3229__A _3232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6583_ _6583_/A _3300_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_3795_ _5484_/A vssd1 vssd1 vccd1 vccd1 _5349_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5534_ _5603_/A _5603_/B _5533_/Y vssd1 vssd1 vccd1 vccd1 _5598_/B sky130_fd_sc_hd__a21o_1
X_5465_ _6278_/Q _5465_/B _5484_/C vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__and3_1
X_4416_ _4266_/A _4430_/B _4392_/C vssd1 vssd1 vccd1 vccd1 _4417_/B sky130_fd_sc_hd__a21oi_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5396_ _5396_/A _5425_/A vssd1 vssd1 vccd1 vccd1 _5397_/B sky130_fd_sc_hd__or2_1
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4347_ _4348_/A _4348_/B vssd1 vssd1 vccd1 vccd1 _4369_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4278_ _4279_/B vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__buf_2
X_3229_ _3232_/A vssd1 vssd1 vccd1 vccd1 _3229_/Y sky130_fd_sc_hd__inv_2
X_6017_ _6026_/A _6017_/B vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__and2_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4507__B _4621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5619__A _5619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5502__A2 _5485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3580_ _3580_/A _4898_/B _3580_/C vssd1 vssd1 vccd1 vccd1 _3580_/Y sky130_fd_sc_hd__nor3_1
X_5250_ _5251_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__nand2_1
X_4201_ _4202_/B _4201_/B vssd1 vssd1 vccd1 vccd1 _4203_/A sky130_fd_sc_hd__and2b_1
XFILLER_5_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5181_ _5174_/A _5180_/X _4062_/A _4961_/B vssd1 vssd1 vccd1 vccd1 _5183_/C sky130_fd_sc_hd__o211ai_4
X_4132_ _4137_/A _4137_/B vssd1 vssd1 vccd1 vccd1 _4138_/C sky130_fd_sc_hd__xor2_1
XFILLER_68_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4063_ _5109_/A _4063_/B _4063_/C vssd1 vssd1 vccd1 vccd1 _4063_/X sky130_fd_sc_hd__and3_1
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4965_ _4972_/B _4972_/A vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4232__A2 _4235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3916_ _3916_/A _3916_/B _3916_/C vssd1 vssd1 vccd1 vccd1 _3917_/B sky130_fd_sc_hd__nand3_1
X_4896_ _3505_/A _4764_/A _4864_/C _3631_/A vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__a22oi_1
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3847_ _5231_/B vssd1 vssd1 vccd1 vccd1 _5195_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _3778_/A _3778_/B vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__nor2_1
X_6566_ _6566_/A _3281_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_5517_ _5648_/A _5641_/B vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__or2_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6497_ _6497_/A _3199_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
X_5448_ _5448_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__xor2_1
X_5379_ _5379_/A _5379_/B vssd1 vssd1 vccd1 vccd1 _5537_/B sky130_fd_sc_hd__xor2_2
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4759__B1 _4796_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6509__28 vssd1 vssd1 vccd1 vccd1 _6509__28/HI _6509_/A sky130_fd_sc_hd__conb_1
XFILLER_8_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3982__A1 _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3332__A _5605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4750_ _3520_/B _4879_/D _4787_/C _3494_/A vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__a22o_1
X_4681_ _4682_/B _4682_/C _4682_/A vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__a21o_1
X_3701_ _3763_/A _3700_/B _3739_/A _3700_/D vssd1 vssd1 vccd1 vccd1 _3702_/C sky130_fd_sc_hd__a22o_1
X_3632_ _3632_/A _5325_/C _3632_/C vssd1 vssd1 vccd1 vccd1 _3632_/X sky130_fd_sc_hd__and3_1
X_6351_ _6359_/CLK _6351_/D vssd1 vssd1 vccd1 vccd1 _6351_/Q sky130_fd_sc_hd__dfxtp_1
X_6523__42 vssd1 vssd1 vccd1 vccd1 _6523__42/HI _6523_/A sky130_fd_sc_hd__conb_1
X_5302_ _5302_/A _5302_/B vssd1 vssd1 vccd1 vccd1 _5339_/B sky130_fd_sc_hd__xnor2_1
X_3563_ _3564_/A _3563_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3583_/A sky130_fd_sc_hd__nand3_1
X_3494_ _3494_/A _3652_/B _3652_/C vssd1 vssd1 vccd1 vccd1 _3495_/B sky130_fd_sc_hd__and3_1
X_6282_ _6345_/CLK _6282_/D vssd1 vssd1 vccd1 vccd1 _6282_/Q sky130_fd_sc_hd__dfxtp_1
X_5233_ _4079_/A _5355_/B _5256_/A _5231_/X vssd1 vssd1 vccd1 vccd1 _5235_/A sky130_fd_sc_hd__a31oi_2
X_5164_ _5382_/C vssd1 vssd1 vccd1 vccd1 _5471_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4115_ _4115_/A _4367_/B _4115_/C vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__and3_1
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5095_ _5070_/B _5091_/Y _5094_/X vssd1 vssd1 vccd1 vccd1 _5123_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3242__A _3245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4046_ _5426_/A vssd1 vssd1 vccd1 vccd1 _5358_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5650__A1 _5511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _5993_/A _5988_/X _5996_/Y _5945_/X vssd1 vssd1 vccd1 vccd1 _6295_/D sky130_fd_sc_hd__o211a_1
X_4948_ _4960_/A _4961_/B _4948_/C vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__and3_1
X_4879_ _4879_/A _4879_/B _4879_/C _4879_/D vssd1 vssd1 vccd1 vccd1 _4897_/A sky130_fd_sc_hd__and4_1
XFILLER_20_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6549_ _6549_/A _3257_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5351__B _5382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_96 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3997__A _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _6098_/A vssd1 vssd1 vccd1 vccd1 _6073_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5851_ _6384_/Q _6283_/Q vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__and2_1
XANTENNA__6092__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4802_ _4802_/A _4802_/B vssd1 vssd1 vccd1 vccd1 _4823_/B sky130_fd_sc_hd__xnor2_1
X_5782_ _6374_/Q _5781_/X _5776_/Y _6375_/Q vssd1 vssd1 vccd1 vccd1 _5782_/X sky130_fd_sc_hd__o22a_1
X_4733_ _4733_/A _4733_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__and3_1
XFILLER_21_248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4664_ _4664_/A _4714_/B _4846_/B vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__and3_1
XANTENNA__3237__A _3239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4595_ _4595_/A _4595_/B vssd1 vssd1 vccd1 vccd1 _4595_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4340__B _4340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3615_ _3615_/A _3615_/B vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__xnor2_1
X_3546_ _3543_/A _3543_/C _3543_/B vssd1 vssd1 vccd1 vccd1 _3621_/B sky130_fd_sc_hd__a21oi_1
X_6334_ _6335_/CLK _6334_/D vssd1 vssd1 vccd1 vccd1 _6334_/Q sky130_fd_sc_hd__dfxtp_1
X_6265_ _6380_/Q _6261_/B _6264_/Y vssd1 vssd1 vccd1 vccd1 _6380_/D sky130_fd_sc_hd__o21a_1
X_5216_ _5198_/A _5215_/X _4323_/A _5236_/B vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__o211a_1
X_3477_ _3696_/A _3652_/B _3652_/C _3477_/D vssd1 vssd1 vccd1 vccd1 _3477_/X sky130_fd_sc_hd__and4_1
XANTENNA__5171__B _5196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6196_ _6196_/A vssd1 vssd1 vccd1 vccd1 _6355_/D sky130_fd_sc_hd__clkbuf_1
X_5147_ _5141_/A _5141_/B _5141_/C vssd1 vssd1 vccd1 vccd1 _5148_/D sky130_fd_sc_hd__a21o_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5078_ _5078_/A _5078_/B _5076_/X vssd1 vssd1 vccd1 vccd1 _5114_/A sky130_fd_sc_hd__or3b_1
X_4029_ _3981_/B _4075_/A _4028_/X vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__o21ai_1
XFILLER_72_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5627__A _5627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4250__B _4250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4380_ _4380_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4384_/B sky130_fd_sc_hd__xor2_1
X_3400_ _3449_/A vssd1 vssd1 vccd1 vccd1 _3400_/X sky130_fd_sc_hd__clkbuf_2
X_3331_ _4548_/A vssd1 vssd1 vccd1 vccd1 _5605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3263_/A vssd1 vssd1 vccd1 vccd1 _3262_/Y sky130_fd_sc_hd__inv_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6050_/A _6051_/A vssd1 vssd1 vccd1 vccd1 _6050_/X sky130_fd_sc_hd__or2b_1
X_5001_ _5001_/A _5145_/B vssd1 vssd1 vccd1 vccd1 _5004_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3193_ _3195_/A vssd1 vssd1 vccd1 vccd1 _3193_/Y sky130_fd_sc_hd__inv_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5903_ _5902_/A _5902_/B _5868_/A vssd1 vssd1 vccd1 vccd1 _5903_/Y sky130_fd_sc_hd__o21ai_1
X_5834_ _6377_/Q _6376_/Q _5834_/C vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__or3_1
X_5765_ input8/X vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__buf_2
X_4716_ _3377_/A _4714_/X _4715_/X vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__a21bo_1
X_5696_ _3396_/Y _4627_/Y _5684_/X _5687_/X _5695_/X vssd1 vssd1 vccd1 vccd1 _5696_/X
+ sky130_fd_sc_hd__a221o_1
X_4647_ _3377_/A _4693_/A _4694_/C vssd1 vssd1 vccd1 vccd1 _4647_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4578_ _5714_/A _4585_/B _4577_/X vssd1 vssd1 vccd1 vccd1 _4578_/Y sky130_fd_sc_hd__a21oi_1
X_6317_ _6384_/CLK _6317_/D vssd1 vssd1 vccd1 vccd1 _6317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3529_ _3529_/A _3529_/B vssd1 vssd1 vccd1 vccd1 _3532_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6248_ _6374_/Q _6373_/Q _6248_/C vssd1 vssd1 vccd1 vccd1 _6249_/B sky130_fd_sc_hd__and3_1
X_6179_ _6348_/Q _6197_/B vssd1 vssd1 vccd1 vccd1 _6180_/A sky130_fd_sc_hd__and2_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4335__A1 _4334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3880_ _3961_/B _3870_/A _3879_/X vssd1 vssd1 vccd1 vccd1 _3965_/B sky130_fd_sc_hd__o21ba_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6565__81 vssd1 vssd1 vccd1 vccd1 _6565__81/HI _6565_/A sky130_fd_sc_hd__conb_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _5550_/A _5550_/B _5550_/C vssd1 vssd1 vccd1 vccd1 _5550_/X sky130_fd_sc_hd__and3_1
X_4501_ _4501_/A _4501_/B vssd1 vssd1 vccd1 vccd1 _4502_/C sky130_fd_sc_hd__or2_1
X_5481_ _5531_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5606_/A sky130_fd_sc_hd__xor2_1
X_4432_ _4411_/A _4429_/Y _4431_/X vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__o21a_1
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4363_ _5349_/A _4153_/C _4372_/A _4361_/X vssd1 vssd1 vccd1 vccd1 _4366_/A sky130_fd_sc_hd__a31o_1
X_3314_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3314_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4294_ _4294_/A _4294_/B vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__nor2_2
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _6102_/A vssd1 vssd1 vccd1 vccd1 _6319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3245_/A vssd1 vssd1 vccd1 vccd1 _3245_/Y sky130_fd_sc_hd__inv_2
X_6033_ _6046_/B vssd1 vssd1 vccd1 vccd1 _6060_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3250__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_298 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5817_ _5813_/X _4627_/Y _5684_/X _5814_/X _5816_/X vssd1 vssd1 vccd1 vccd1 _5817_/X
+ sky130_fd_sc_hd__a221o_1
X_5748_ _5671_/Y _5674_/Y _5677_/Y vssd1 vssd1 vccd1 vccd1 _5749_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_448 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5679_ _5679_/A vssd1 vssd1 vccd1 vccd1 _5719_/A sky130_fd_sc_hd__inv_2
XFILLER_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5293__A2 _5485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5640__A _5646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5348__A3 _5471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4556__A1 _5698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4166__A _5355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4981_ _4981_/A _4964_/B vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__or2b_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _4488_/A _3932_/B vssd1 vssd1 vccd1 vccd1 _3934_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ _3885_/C _3863_/B vssd1 vssd1 vccd1 vccd1 _3864_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__4547__A1 _4546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5602_ _5737_/A _5652_/A vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__xnor2_1
X_6582_ _6582_/A _3299_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3794_ _6276_/Q vssd1 vssd1 vccd1 vccd1 _5484_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5533_ _5533_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5533_/Y sky130_fd_sc_hd__nor2_1
X_5464_ _5464_/A _5464_/B vssd1 vssd1 vccd1 vccd1 _5478_/A sky130_fd_sc_hd__xor2_1
XFILLER_99_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4415_ _4415_/A vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__inv_2
X_5395_ _5396_/A _5425_/A vssd1 vssd1 vccd1 vccd1 _5397_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5444__B _5444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4346_ _4346_/A _4346_/B vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3245__A _3245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4277_ _4312_/A _5450_/C vssd1 vssd1 vccd1 vccd1 _4279_/B sky130_fd_sc_hd__and2_1
X_6016_ _6016_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__or2_1
X_3228_ _3232_/A vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5027__A2 _5013_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6293__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5974__B1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5726__B1 _5737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4200_ _4198_/A _4198_/B _4240_/A vssd1 vssd1 vccd1 vccd1 _4201_/B sky130_fd_sc_hd__o21ai_1
XFILLER_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _5174_/A _5174_/B _5180_/C _5180_/D vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__and4bb_1
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4131_ _5404_/A _4131_/B vssd1 vssd1 vccd1 vccd1 _4137_/B sky130_fd_sc_hd__and2_1
XFILLER_68_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4062_ _4062_/A vssd1 vssd1 vccd1 vccd1 _5109_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4964_ _4981_/A _4964_/B vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__xnor2_1
X_3915_ _3916_/A _3916_/B _3916_/C vssd1 vssd1 vccd1 vccd1 _3934_/A sky130_fd_sc_hd__a21o_1
X_4895_ _4895_/A _4895_/B vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3846_ _5312_/A vssd1 vssd1 vccd1 vccd1 _5231_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3777_ _3777_/A _3777_/B vssd1 vssd1 vccd1 vccd1 _3778_/B sky130_fd_sc_hd__and2_1
X_6565_ _6565_/A _3280_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
X_5516_ _5516_/A _5516_/B vssd1 vssd1 vccd1 vccd1 _5641_/B sky130_fd_sc_hd__or2_1
X_6496_ _6496_/A _3198_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
X_5447_ _5447_/A _5447_/B vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5496__A2 _5489_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5378_ _5539_/B _5378_/B vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__xnor2_4
XFILLER_87_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4329_ _4329_/A _4329_/B vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__xor2_4
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4759__B2 _3601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__B _5444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3982__A2 _4168_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5184__A1 _4059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5365__A _5505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_187 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _3763_/A _3700_/B _3739_/A _3700_/D vssd1 vssd1 vccd1 vccd1 _3739_/B sky130_fd_sc_hd__nand4_1
X_4680_ _4680_/A _4680_/B vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5175__B2 _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ _3631_/A _5450_/C vssd1 vssd1 vccd1 vccd1 _5325_/C sky130_fd_sc_hd__nand2_1
X_6350_ _6357_/CLK _6350_/D vssd1 vssd1 vccd1 vccd1 _6350_/Q sky130_fd_sc_hd__dfxtp_1
X_3562_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3563_/C sky130_fd_sc_hd__xor2_1
X_5301_ _5301_/A _5301_/B vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__xor2_1
X_3493_ _3690_/A _3696_/B vssd1 vssd1 vccd1 vccd1 _3495_/A sky130_fd_sc_hd__nand2_1
X_6281_ _6359_/CLK _6281_/D vssd1 vssd1 vccd1 vccd1 _6281_/Q sky130_fd_sc_hd__dfxtp_1
X_5232_ _5196_/C _5230_/X _5231_/X vssd1 vssd1 vccd1 vccd1 _5256_/A sky130_fd_sc_hd__o21ba_1
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _5161_/A _5161_/B _4909_/X vssd1 vssd1 vccd1 vccd1 _5382_/C sky130_fd_sc_hd__o21bai_2
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4114_ _4114_/A _4153_/B vssd1 vssd1 vccd1 vccd1 _4115_/C sky130_fd_sc_hd__xor2_1
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5094_ _5091_/A _5388_/B _5130_/B vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__a21o_1
X_4045_ _5489_/A vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _5994_/X _5995_/Y _6057_/A vssd1 vssd1 vccd1 vccd1 _5996_/Y sky130_fd_sc_hd__o21ai_1
X_4947_ _4947_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4948_/C sky130_fd_sc_hd__xor2_1
XANTENNA__4073__B _4365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4878_ _4842_/A _4879_/C _4877_/D _3645_/B vssd1 vssd1 vccd1 vccd1 _4881_/B sky130_fd_sc_hd__a22o_1
X_3829_ _3826_/B _3829_/B vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6548_ _6548_/A _3260_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_552 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_680 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3608__A _4882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4904__B2 _4726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5632__A2 _5630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5850_ _6383_/Q _5818_/Y _5823_/X _5849_/X _6259_/A vssd1 vssd1 vccd1 vccd1 _6536_/A
+ sky130_fd_sc_hd__a221oi_4
X_4801_ _4801_/A _4801_/B vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__or2_1
X_5781_ _5698_/A _5778_/X _5780_/X _5706_/X vssd1 vssd1 vccd1 vccd1 _5781_/X sky130_fd_sc_hd__o2bb2a_1
X_4732_ _4732_/A _4755_/A vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__xnor2_4
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__4621__B _4621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _3634_/B _3614_/B vssd1 vssd1 vccd1 vccd1 _3614_/Y sky130_fd_sc_hd__nor2_1
X_4594_ _4370_/B _4606_/B _4592_/B _5740_/A vssd1 vssd1 vccd1 vccd1 _4594_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3545_ _3640_/B _3545_/B vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__xnor2_1
X_6333_ _6359_/CLK _6333_/D vssd1 vssd1 vccd1 vccd1 _6333_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5733__A _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3476_ _3465_/B _3465_/C _3465_/A vssd1 vssd1 vccd1 vccd1 _3476_/Y sky130_fd_sc_hd__a21boi_1
X_6264_ _6267_/A _6269_/C vssd1 vssd1 vccd1 vccd1 _6264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5215_ _5215_/A _5215_/B _5215_/C vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__and3_1
XANTENNA__3253__A _3257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6195_ _6354_/Q _6197_/B vssd1 vssd1 vccd1 vccd1 _6196_/A sky130_fd_sc_hd__and2_1
XFILLER_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5146_ _5183_/A _5109_/B _5151_/A _5145_/D vssd1 vssd1 vccd1 vccd1 _5148_/C sky130_fd_sc_hd__a22o_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5077_ _5078_/A _5078_/B _5076_/X vssd1 vssd1 vccd1 vccd1 _5114_/C sky130_fd_sc_hd__o21bai_1
XFILLER_29_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4028_ _5130_/A _4323_/B _4367_/B _5129_/A vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5979_ _5979_/A vssd1 vssd1 vccd1 vccd1 _6292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3428__A _6040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3873__B2 _5001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3338__A _4933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5040__D_N _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _4974_/A vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5634_/A _5000_/B vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__nand2_1
X_3261_ _3263_/A vssd1 vssd1 vccd1 vccd1 _3261_/Y sky130_fd_sc_hd__inv_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3195_/A vssd1 vssd1 vccd1 vccd1 _3192_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5902_ _5902_/A _5902_/B vssd1 vssd1 vccd1 vccd1 _5902_/X sky130_fd_sc_hd__and2_1
XFILLER_62_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5833_ _6376_/Q _5834_/C _6258_/B vssd1 vssd1 vccd1 vccd1 _5833_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4632__A _4769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5764_ _5754_/X _5762_/X _5763_/X vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__a21o_1
X_4715_ _4714_/A _4714_/B _4785_/C _4645_/A vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3248__A _3251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5695_ _5613_/A _5699_/B _5694_/X vssd1 vssd1 vccd1 vccd1 _5695_/X sky130_fd_sc_hd__a21o_1
X_4646_ _4714_/A _4692_/B vssd1 vssd1 vccd1 vccd1 _4694_/C sky130_fd_sc_hd__nand2_1
XFILLER_30_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4577_ _4577_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _4577_/X sky130_fd_sc_hd__and2_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _6369_/CLK _6316_/D vssd1 vssd1 vccd1 vccd1 _6316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3528_ _4846_/A _3692_/B vssd1 vssd1 vccd1 vccd1 _3540_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6247_ _6373_/Q _6248_/C _6246_/Y vssd1 vssd1 vccd1 vccd1 _6373_/D sky130_fd_sc_hd__o21a_1
X_3459_ _4842_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3464_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6178_ _6178_/A vssd1 vssd1 vccd1 vccd1 _6197_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5129_ _5129_/A _5243_/B vssd1 vssd1 vccd1 vccd1 _5129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5092__B _5355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4099__A1 _4138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4717__A _5966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5707__A1_N _5906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5267__B _5267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4500_ _4141_/B _4141_/C _4141_/A vssd1 vssd1 vccd1 vccd1 _4501_/B sky130_fd_sc_hd__a21oi_1
X_5480_ _5478_/A _5478_/B _5479_/X vssd1 vssd1 vccd1 vccd1 _5531_/B sky130_fd_sc_hd__o21a_1
X_4431_ _5510_/A _4153_/C _4445_/A vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__a21bo_1
XFILLER_6_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6580__96 vssd1 vssd1 vccd1 vccd1 _6580__96/HI _6580_/A sky130_fd_sc_hd__conb_1
XFILLER_6_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4362_ _4332_/B _4359_/Y _4361_/X vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__a21oi_1
XFILLER_112_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3313_ _3313_/A vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__buf_6
X_4293_ _4296_/A _4296_/B vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__and2b_1
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _6318_/Q _6107_/B vssd1 vssd1 vccd1 vccd1 _6102_/A sky130_fd_sc_hd__and2_1
XFILLER_112_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3244_ _3245_/A vssd1 vssd1 vccd1 vccd1 _3244_/Y sky130_fd_sc_hd__inv_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6042_/A _6032_/B vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__and2_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5816_ _5613_/A _5819_/B _5694_/X vssd1 vssd1 vccd1 vccd1 _5816_/X sky130_fd_sc_hd__a21o_1
X_5747_ _5747_/A _5747_/B vssd1 vssd1 vccd1 vccd1 _5747_/X sky130_fd_sc_hd__and2_1
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _5671_/Y _5674_/Y _5749_/A _5677_/Y vssd1 vssd1 vccd1 vccd1 _5678_/X sky130_fd_sc_hd__o211a_1
X_4629_ _4726_/B vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_116_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4166__B _4166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _4988_/B _4980_/B vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__or2_1
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5278__A _5278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3931_ _3931_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _3932_/B sky130_fd_sc_hd__or2_1
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3862_ _4925_/A _4131_/B vssd1 vssd1 vccd1 vccd1 _3863_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6581_ _6581_/A _3298_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
XANTENNA__4547__A2 _4546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5601_ _5601_/A _5601_/B vssd1 vssd1 vccd1 vccd1 _5601_/Y sky130_fd_sc_hd__nand2_1
X_3793_ _3793_/A _3793_/B vssd1 vssd1 vccd1 vccd1 _3939_/A sky130_fd_sc_hd__xnor2_1
X_5532_ _5606_/A _5606_/B _5531_/Y vssd1 vssd1 vccd1 vccd1 _5603_/B sky130_fd_sc_hd__a21o_1
X_5463_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5464_/B sky130_fd_sc_hd__xnor2_1
X_4414_ _5314_/A _4153_/C _4435_/A _4413_/X vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__a31o_1
XANTENNA__5444__C _5444_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5394_ _5394_/A _5394_/B _5484_/C vssd1 vssd1 vccd1 vccd1 _5425_/A sky130_fd_sc_hd__and3_1
X_4345_ _4374_/A _4374_/B vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__and2_1
XFILLER_98_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4276_ _4276_/A _4276_/B vssd1 vssd1 vccd1 vccd1 _4284_/B sky130_fd_sc_hd__xor2_1
X_3227_ _3227_/A vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__buf_8
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3261__A _3263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6015_ _6016_/A _6031_/B vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5101__D_N _5059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_244 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5974__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5264__C _5267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6550__66 vssd1 vssd1 vccd1 vccd1 _6550__66/HI _6550_/A sky130_fd_sc_hd__conb_1
X_4130_ _5276_/A vssd1 vssd1 vccd1 vccd1 _5404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4061_ _4138_/A vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ _4975_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _4964_/B sky130_fd_sc_hd__xor2_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3914_ _3931_/A _3913_/X vssd1 vssd1 vccd1 vccd1 _3916_/C sky130_fd_sc_hd__or2b_1
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4894_ _4894_/A _4894_/B _4894_/C vssd1 vssd1 vccd1 vccd1 _4895_/B sky130_fd_sc_hd__and3_1
X_3845_ _4331_/A vssd1 vssd1 vccd1 vccd1 _5312_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3776_ _3777_/A _3777_/B vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__nor2_1
X_6564_ _6564_/A _3279_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_5515_ _5514_/B _5514_/C _5514_/A vssd1 vssd1 vccd1 vccd1 _5516_/B sky130_fd_sc_hd__a21oi_1
X_6495_ _6495_/A _3197_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
XFILLER_105_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3256__A _3257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5446_ _5463_/A _5463_/B vssd1 vssd1 vccd1 vccd1 _5447_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5377_ _5379_/A _5379_/B _5376_/X vssd1 vssd1 vccd1 vccd1 _5378_/B sky130_fd_sc_hd__a21oi_2
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4328_ _4465_/B _4328_/B vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__xnor2_4
X_4259_ _4469_/A _4469_/B vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__xor2_4
XANTENNA_input1_A active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5349__C _5444_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5646__A _5646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__B _4769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ _4820_/B vssd1 vssd1 vccd1 vccd1 _5450_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3561_ _3560_/A _3560_/B _3560_/C vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__a21o_1
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5300_ _5300_/A _5300_/B vssd1 vssd1 vccd1 vccd1 _5339_/A sky130_fd_sc_hd__xor2_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6280_ _6359_/CLK _6280_/D vssd1 vssd1 vccd1 vccd1 _6280_/Q sky130_fd_sc_hd__dfxtp_1
X_3492_ _3492_/A vssd1 vssd1 vccd1 vccd1 _3696_/B sky130_fd_sc_hd__clkbuf_2
X_5231_ _5231_/A _5231_/B _5273_/B _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__and4_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5162_ _5382_/B vssd1 vssd1 vccd1 vccd1 _5471_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _5166_/A _5231_/D vssd1 vssd1 vccd1 vccd1 _5130_/B sky130_fd_sc_hd__and2_1
X_4113_ _4194_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4153_/B sky130_fd_sc_hd__and2_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4044_ _5510_/A vssd1 vssd1 vccd1 vccd1 _5489_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6283__CLK _6384_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5995_ _5995_/A _5995_/B vssd1 vssd1 vccd1 vccd1 _5995_/Y sky130_fd_sc_hd__nor2_1
X_4946_ _5218_/D vssd1 vssd1 vccd1 vccd1 _4961_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4877_ _4877_/A _4877_/B _4877_/C _4877_/D vssd1 vssd1 vccd1 vccd1 _4881_/A sky130_fd_sc_hd__nand4_1
X_3828_ _3825_/A _3825_/B _3827_/Y _3822_/X vssd1 vssd1 vccd1 vccd1 _3828_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4370__A _5246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6547_ _6547_/A _3262_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
X_3759_ _3742_/B _3759_/B vssd1 vssd1 vccd1 vccd1 _3759_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6514__33 vssd1 vssd1 vccd1 vccd1 _6514__33/HI _6514_/A sky130_fd_sc_hd__conb_1
X_5429_ _5429_/A _5429_/B vssd1 vssd1 vccd1 vccd1 _5448_/B sky130_fd_sc_hd__xnor2_1
XFILLER_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4529__B _4577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_114 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_64 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4264__B _4412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4904__A2 _4898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4668__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4800_ _4818_/A _4800_/B vssd1 vssd1 vccd1 vccd1 _4801_/B sky130_fd_sc_hd__nor2_1
X_5780_ _5690_/A _5703_/Y _5815_/B _5702_/Y vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__o22a_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4731_/A _4731_/B _4764_/A _4796_/D vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__and4_2
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662_ _4662_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__nor2_1
X_3613_ _3633_/A _3613_/B vssd1 vssd1 vccd1 vccd1 _3614_/B sky130_fd_sc_hd__nand2_1
X_4593_ _4593_/A _4593_/B vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__xor2_2
X_3544_ _3544_/A _3621_/A vssd1 vssd1 vccd1 vccd1 _3545_/B sky130_fd_sc_hd__nor2_1
X_6332_ _6345_/CLK _6332_/D vssd1 vssd1 vccd1 vccd1 _6332_/Q sky130_fd_sc_hd__dfxtp_1
X_3475_ _3536_/A _3536_/B _3536_/C vssd1 vssd1 vccd1 vccd1 _3475_/Y sky130_fd_sc_hd__nand3_1
X_6263_ _6380_/Q _6379_/Q _6263_/C vssd1 vssd1 vccd1 vccd1 _6269_/C sky130_fd_sc_hd__and3_1
X_5214_ _5214_/A _5214_/B _5213_/X vssd1 vssd1 vccd1 vccd1 _5221_/A sky130_fd_sc_hd__nor3b_2
X_6194_ _6194_/A vssd1 vssd1 vccd1 vccd1 _6354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5145_ _5183_/A _5145_/B _5151_/A _5145_/D vssd1 vssd1 vccd1 vccd1 _5151_/B sky130_fd_sc_hd__nand4_1
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5074_/A _5074_/B _5107_/A vssd1 vssd1 vccd1 vccd1 _5076_/X sky130_fd_sc_hd__a21bo_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _4376_/B vssd1 vssd1 vccd1 vccd1 _4367_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _6350_/Q _5980_/B vssd1 vssd1 vccd1 vccd1 _5979_/A sky130_fd_sc_hd__and2_1
X_4929_ _4929_/A _5180_/D vssd1 vssd1 vccd1 vccd1 _4947_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5311__A2 _5444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6272__B1 _6218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3260_ _3263_/A vssd1 vssd1 vccd1 vccd1 _3260_/Y sky130_fd_sc_hd__inv_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3191_ _3195_/A vssd1 vssd1 vccd1 vccd1 _3191_/Y sky130_fd_sc_hd__inv_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5901_ _5901_/A _5906_/B vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__xnor2_1
XFILLER_81_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _6377_/Q vssd1 vssd1 vccd1 vccd1 _6258_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5763_ _6365_/Q _5761_/X _5707_/X _6366_/Q vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__a22o_1
X_4714_ _4714_/A _4714_/B _4785_/C vssd1 vssd1 vccd1 vccd1 _4714_/X sky130_fd_sc_hd__and3_1
X_5694_ _5841_/B vssd1 vssd1 vccd1 vccd1 _5694_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4645_ _4645_/A _4645_/B _4675_/C _4692_/B vssd1 vssd1 vccd1 vccd1 _4645_/Y sky130_fd_sc_hd__nand4_2
XFILLER_30_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4576_ _4577_/A _4577_/B vssd1 vssd1 vccd1 vccd1 _4585_/B sky130_fd_sc_hd__xor2_1
X_6315_ _6384_/CLK _6315_/D vssd1 vssd1 vccd1 vccd1 _6315_/Q sky130_fd_sc_hd__dfxtp_1
X_3527_ _3527_/A _3560_/A vssd1 vssd1 vccd1 vccd1 _3565_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3264__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6246_ _6267_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6246_/Y sky130_fd_sc_hd__nor2_1
X_3458_ _3458_/A _3653_/C vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__and2_1
XFILLER_76_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6177_ _6177_/A vssd1 vssd1 vccd1 vccd1 _6348_/D sky130_fd_sc_hd__clkbuf_1
X_3389_ _5813_/B vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__clkbuf_2
X_5128_ _5274_/D vssd1 vssd1 vccd1 vccd1 _5243_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5059_/A _5059_/B _5059_/C vssd1 vssd1 vccd1 vccd1 _5062_/A sky130_fd_sc_hd__and3_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4099__A2 _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4717__B _4814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ _5485_/A _4430_/B vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4361_ _5411_/A _4361_/B _4361_/C vssd1 vssd1 vccd1 vccd1 _4361_/X sky130_fd_sc_hd__and3_1
XFILLER_6_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6100_ _6100_/A vssd1 vssd1 vccd1 vccd1 _6318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4292_ _4292_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4296_/B sky130_fd_sc_hd__xnor2_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _3312_/A vssd1 vssd1 vccd1 vccd1 _3312_/Y sky130_fd_sc_hd__inv_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3245_/A vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__inv_2
X_6031_ _6300_/Q _6031_/B vssd1 vssd1 vccd1 vccd1 _6032_/B sky130_fd_sc_hd__or2_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5039__A1 _5001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5815_ _5815_/A _5815_/B vssd1 vssd1 vccd1 vccd1 _5819_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3259__A _3263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6556__72 vssd1 vssd1 vccd1 vccd1 _6556__72/HI _6556_/A sky130_fd_sc_hd__conb_1
X_5746_ _5746_/A _5746_/B _5746_/C vssd1 vssd1 vccd1 vccd1 _5747_/B sky130_fd_sc_hd__nand3_1
XFILLER_41_28 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5677_ _5677_/A _5677_/B vssd1 vssd1 vccd1 vccd1 _5677_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4628_ _4796_/D vssd1 vssd1 vccd1 vccd1 _4726_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_104_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4559_ _4559_/A _4559_/B vssd1 vssd1 vccd1 vccd1 _4561_/B sky130_fd_sc_hd__and2_1
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4818__A _4818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6229_ _6366_/Q _6225_/B _6228_/Y vssd1 vssd1 vccd1 vccd1 _6366_/D sky130_fd_sc_hd__o21a_1
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _3931_/A _3931_/B vssd1 vssd1 vccd1 vccd1 _4488_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5278__B _5278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3861_ _5007_/A vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3792_ _3792_/A _3792_/B vssd1 vssd1 vccd1 vccd1 _3793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5600_ _5727_/A _5644_/A vssd1 vssd1 vccd1 vccd1 _5601_/B sky130_fd_sc_hd__nand2_1
X_6580_ _6580_/A _3296_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5531_ _5531_/A _5531_/B vssd1 vssd1 vccd1 vccd1 _5531_/Y sky130_fd_sc_hd__nor2_1
X_5462_ _5462_/A _5462_/B vssd1 vssd1 vccd1 vccd1 _5531_/A sky130_fd_sc_hd__xnor2_1
X_4413_ _4418_/A _4418_/B vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__and2b_1
X_5393_ _5393_/A _5393_/B vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__xnor2_1
X_4344_ _4344_/A _4344_/B vssd1 vssd1 vccd1 vccd1 _4374_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4275_ _4275_/A _4275_/B vssd1 vssd1 vccd1 vccd1 _4276_/B sky130_fd_sc_hd__nor2_1
X_6014_ _6297_/Q _5988_/X _6012_/Y _6013_/X vssd1 vssd1 vccd1 vccd1 _6297_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3226_ _3226_/A vssd1 vssd1 vccd1 vccd1 _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _6362_/Q vssd1 vssd1 vccd1 vccd1 _5729_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5098__B _5099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3362__A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4060_ _5183_/A vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _4974_/A _5013_/B vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _3913_/A _3913_/B _3911_/X vssd1 vssd1 vccd1 vccd1 _3913_/X sky130_fd_sc_hd__or3b_1
X_4893_ _4891_/A _4890_/C _4890_/B vssd1 vssd1 vccd1 vccd1 _4908_/B sky130_fd_sc_hd__a21o_1
X_3844_ _5410_/A vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3775_ _3804_/A _3804_/B vssd1 vssd1 vccd1 vccd1 _3777_/B sky130_fd_sc_hd__xnor2_1
X_6563_ _6563_/A _3278_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
XFILLER_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5514_ _5514_/A _5514_/B _5514_/C vssd1 vssd1 vccd1 vccd1 _5516_/A sky130_fd_sc_hd__and3_1
X_6494_ _6494_/A _3195_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5445_ _5445_/A _5445_/B vssd1 vssd1 vccd1 vccd1 _5463_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5376_ _5375_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5376_/X sky130_fd_sc_hd__and2b_1
XANTENNA__5471__B _5471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3272__A _3276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4327_ _4322_/A _4322_/B _4326_/X vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__o21ba_2
X_4258_ _4260_/A _4260_/B _4257_/Y vssd1 vssd1 vccd1 vccd1 _4469_/B sky130_fd_sc_hd__a21o_2
XFILLER_47_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3209_ _3227_/A vssd1 vssd1 vccd1 vccd1 _3214_/A sky130_fd_sc_hd__buf_6
XFILLER_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4189_ _4189_/A _4189_/B vssd1 vssd1 vccd1 vccd1 _4202_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5405__A1 _5355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5381__B _5486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3357__A _6291_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3560_ _3560_/A _3560_/B _3560_/C vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__nand3_1
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230_ _5230_/A _5231_/D vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__and2_1
X_3491_ _4877_/B _3692_/B vssd1 vssd1 vccd1 vccd1 _3496_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5161_ _5161_/A _5161_/B _4909_/X vssd1 vssd1 vccd1 vccd1 _5382_/B sky130_fd_sc_hd__or3b_2
XFILLER_110_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5092_ _5158_/A _5355_/B vssd1 vssd1 vccd1 vccd1 _5123_/A sky130_fd_sc_hd__nand2_1
X_4112_ _4110_/X _4111_/X _4072_/C vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__o21a_2
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4043_ _6274_/Q vssd1 vssd1 vccd1 vccd1 _5510_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _5995_/A _5995_/B vssd1 vssd1 vccd1 vccd1 _5994_/X sky130_fd_sc_hd__and2_1
X_4945_ _5059_/B vssd1 vssd1 vccd1 vccd1 _5218_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4876_ _4869_/A _4869_/C _4869_/B vssd1 vssd1 vccd1 vccd1 _4889_/C sky130_fd_sc_hd__a21o_1
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3827_ _3484_/A _3503_/B _3764_/B vssd1 vssd1 vccd1 vccd1 _3827_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4370__B _4370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3267__A _3270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3758_ _3758_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3777_/A sky130_fd_sc_hd__nand2_1
X_6546_ _6546_/A _3266_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
X_3689_ _3657_/B _3657_/C _3657_/A vssd1 vssd1 vccd1 vccd1 _3706_/A sky130_fd_sc_hd__a21bo_1
X_5428_ _5449_/A _5449_/B vssd1 vssd1 vccd1 vccd1 _5429_/B sky130_fd_sc_hd__or2_1
XFILLER_114_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5359_ _5359_/A _5359_/B vssd1 vssd1 vccd1 vccd1 _5380_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5657__A _5885_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6000__B _6000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4668__A2 _5685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5617__A1 _5698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4877_/C vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__clkbuf_2
X_4661_ _4660_/B _4689_/A vssd1 vssd1 vccd1 vccd1 _4662_/B sky130_fd_sc_hd__and2b_1
X_3612_ _3632_/A _3632_/C vssd1 vssd1 vccd1 vccd1 _3613_/B sky130_fd_sc_hd__nor2_1
X_4592_ _5740_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _4595_/B sky130_fd_sc_hd__nand2_1
X_6331_ _6345_/CLK _6331_/D vssd1 vssd1 vccd1 vccd1 _6331_/Q sky130_fd_sc_hd__dfxtp_1
X_3543_ _3543_/A _3543_/B _3543_/C vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__and3_1
X_3474_ _3474_/A _3474_/B vssd1 vssd1 vccd1 vccd1 _3536_/C sky130_fd_sc_hd__nor2_1
X_6262_ _6379_/Q _6263_/C _6261_/Y vssd1 vssd1 vccd1 vccd1 _6379_/D sky130_fd_sc_hd__o21a_1
X_5213_ _5242_/A _5242_/B _5212_/A vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__a21o_1
X_6193_ _6353_/Q _6197_/B vssd1 vssd1 vccd1 vccd1 _6194_/A sky130_fd_sc_hd__and2_1
X_5144_ _4053_/A _5038_/B _5136_/A _5142_/Y vssd1 vssd1 vccd1 vccd1 _5145_/D sky130_fd_sc_hd__a211o_1
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5075_ _5075_/A _5075_/B _5075_/C vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__nand3_1
XANTENNA__3550__A _6284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4026_ _4334_/B vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ _5977_/A vssd1 vssd1 vccd1 vccd1 _6291_/D sky130_fd_sc_hd__clkbuf_1
X_4928_ _5278_/B vssd1 vssd1 vccd1 vccd1 _5180_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5196__B _5196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4856_/X _4857_/X _4860_/A _4858_/Y vssd1 vssd1 vccd1 vccd1 _4860_/B sky130_fd_sc_hd__a211oi_2
XANTENNA__3428__C _4707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3725__A _5246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6529_ _6529_/A _3238_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
XFILLER_106_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5311__A3 _5444_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4035__B1 _3987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_354 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3195_/A sky130_fd_sc_hd__buf_8
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5900_ _5892_/B _5895_/B _5899_/Y vssd1 vssd1 vccd1 vccd1 _5902_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__3520__D _5325_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5831_ _5866_/A _5820_/A _5830_/X _5715_/B vssd1 vssd1 vccd1 vccd1 _5834_/C sky130_fd_sc_hd__a22oi_2
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5762_ _6364_/Q _5713_/Y _5761_/X _6365_/Q vssd1 vssd1 vccd1 vccd1 _5762_/X sky130_fd_sc_hd__o22a_1
X_4713_ _4719_/A _4719_/B _4719_/C vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__a21o_1
X_5693_ _5777_/A vssd1 vssd1 vccd1 vccd1 _5841_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4644_ _4644_/A _4645_/A _4693_/A _4692_/B vssd1 vssd1 vccd1 vccd1 _4656_/B sky130_fd_sc_hd__and4_1
X_4575_ _4575_/A _4575_/B vssd1 vssd1 vccd1 vccd1 _4577_/B sky130_fd_sc_hd__nor2_1
X_6314_ _6384_/CLK _6314_/D vssd1 vssd1 vccd1 vccd1 _6314_/Q sky130_fd_sc_hd__dfxtp_1
X_3526_ _3516_/Y _3529_/B _3526_/C vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__nand3b_1
XFILLER_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6245_ _6373_/Q _6248_/C vssd1 vssd1 vccd1 vccd1 _6246_/B sky130_fd_sc_hd__and2_1
XFILLER_103_359 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3457_ _6016_/A _3400_/X _4749_/A _4641_/A vssd1 vssd1 vccd1 vccd1 _3653_/C sky130_fd_sc_hd__o31ai_2
X_6176_ _6347_/Q _6176_/B vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__and2_1
X_3388_ _5779_/A vssd1 vssd1 vccd1 vccd1 _5813_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5127_ _5269_/A _5270_/A vssd1 vssd1 vccd1 vccd1 _5274_/D sky130_fd_sc_hd__and2_1
X_5058_ _5097_/A _5099_/A vssd1 vssd1 vccd1 vccd1 _5059_/C sky130_fd_sc_hd__and2_1
XANTENNA__3280__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _4009_/A _4009_/B vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5000__A _5634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5935__A _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__6296__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3190__A _3321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5756__B1 _4626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_10 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4360_ _5410_/A _4388_/B vssd1 vssd1 vccd1 vccd1 _4361_/C sky130_fd_sc_hd__and2_1
XFILLER_6_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3311_ _3312_/A vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__inv_2
X_4291_ _4270_/B _4272_/B _4270_/A vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__o21ba_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3245_/A vssd1 vssd1 vccd1 vccd1 _3242_/Y sky130_fd_sc_hd__inv_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6300_/Q _6046_/B vssd1 vssd1 vccd1 vccd1 _6042_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4924__A _5099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5814_ _5813_/B _6060_/A _5814_/C vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__and3b_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5755__A _5755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5745_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5867_/A sky130_fd_sc_hd__clkbuf_2
X_5676_ _5676_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _5749_/A sky130_fd_sc_hd__xnor2_1
X_4627_ _5702_/A _5757_/A _4516_/A vssd1 vssd1 vccd1 vccd1 _4627_/Y sky130_fd_sc_hd__o21ai_2
X_6571__87 vssd1 vssd1 vccd1 vccd1 _6571__87/HI _6571_/A sky130_fd_sc_hd__conb_1
XANTENNA__3275__A _3276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4558_ _4558_/A _4558_/B _4566_/A vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__nand3_1
XFILLER_104_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4489_ _4496_/A _4489_/B vssd1 vssd1 vccd1 vccd1 _4490_/B sky130_fd_sc_hd__xor2_4
X_3509_ _3508_/A _3508_/B _3507_/X vssd1 vssd1 vccd1 vccd1 _3509_/X sky130_fd_sc_hd__o21ba_1
X_6228_ _6242_/A _6228_/B vssd1 vssd1 vccd1 vccd1 _6228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3722__B _4235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6334_/Q _6333_/Q _6336_/Q vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__or3_1
XFILLER_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_40 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3860_ _4128_/B vssd1 vssd1 vccd1 vccd1 _4138_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3791_ _3754_/B _3885_/C _3790_/X vssd1 vssd1 vccd1 vccd1 _3792_/B sky130_fd_sc_hd__a21boi_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5530_ _5614_/A _5622_/A _5529_/X vssd1 vssd1 vccd1 vccd1 _5606_/B sky130_fd_sc_hd__o21ai_1
X_5461_ _5533_/A _5533_/B vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__xor2_2
X_4412_ _6274_/Q _4412_/B vssd1 vssd1 vccd1 vccd1 _4418_/B sky130_fd_sc_hd__and2_1
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5392_ _5367_/X _5392_/B vssd1 vssd1 vccd1 vccd1 _5393_/B sky130_fd_sc_hd__and2b_1
X_4343_ _5450_/B _4580_/B _5394_/B vssd1 vssd1 vccd1 vccd1 _4344_/B sky130_fd_sc_hd__a21oi_1
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4274_ _4274_/A _4274_/B vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3225_ _3226_/A vssd1 vssd1 vccd1 vccd1 _3225_/Y sky130_fd_sc_hd__inv_2
X_6013_ _6187_/A vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5469__B _5469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _3994_/A _3994_/B vssd1 vssd1 vccd1 vccd1 _4040_/B sky130_fd_sc_hd__xor2_1
X_5728_ _3396_/Y _5724_/Y _5727_/Y _5687_/X vssd1 vssd1 vccd1 vccd1 _5728_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5659_ _5659_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6334__CLK _6335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4564__A _5627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3434__A1 _5935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_6535__54 vssd1 vssd1 vccd1 vccd1 _6535__54/HI _6535_/A sky130_fd_sc_hd__conb_1
XFILLER_114_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4961_ _4961_/A _4961_/B vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3425__A1 _3387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4892_ _4910_/A _4910_/B _4910_/C vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__a21o_1
X_3912_ _3913_/A _3913_/B _3911_/X vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__o21ba_1
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3843_ _6277_/Q vssd1 vssd1 vccd1 vccd1 _5410_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6562_ _6562_/A _3276_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_3774_ _3774_/A _3774_/B vssd1 vssd1 vccd1 vccd1 _3804_/B sky130_fd_sc_hd__xnor2_1
X_5513_ _5471_/A _5365_/X _5510_/B _4334_/A vssd1 vssd1 vccd1 vccd1 _5514_/C sky130_fd_sc_hd__a22o_1
X_6493_ _6493_/A _3194_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
X_5444_ _5471_/A _5444_/B _5444_/C vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__and3_1
X_6541__57 vssd1 vssd1 vccd1 vccd1 _6541__57/HI _6541_/A sky130_fd_sc_hd__conb_1
XFILLER_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5375_ _5375_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5379_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__5471__C _5471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _4329_/B _4329_/A vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__and2b_1
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4257_ _4257_/A _4257_/B vssd1 vssd1 vccd1 vccd1 _4257_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5102__B2 _5059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3208_ _3208_/A vssd1 vssd1 vccd1 vccd1 _3208_/Y sky130_fd_sc_hd__inv_2
X_4188_ _4188_/A _4188_/B vssd1 vssd1 vccd1 vccd1 _4189_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3728__A _5085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3490_ _3643_/B _3489_/C _3489_/A vssd1 vssd1 vccd1 vccd1 _3497_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _4910_/A _4910_/B _4910_/C vssd1 vssd1 vccd1 vccd1 _5161_/B sky130_fd_sc_hd__a21oi_1
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5091_ _5091_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _5091_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4111_ _3629_/A _3614_/Y _3635_/B vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__a21o_1
X_4042_ _4042_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _4097_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5993_ _5993_/A _6000_/B vssd1 vssd1 vccd1 vccd1 _5995_/B sky130_fd_sc_hd__xor2_1
X_4944_ _4944_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _5059_/B sky130_fd_sc_hd__xnor2_4
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4875_ _4873_/A _4873_/C _4873_/B vssd1 vssd1 vccd1 vccd1 _4910_/B sky130_fd_sc_hd__a21o_1
X_3826_ _3829_/B _3826_/B vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__xnor2_4
X_3757_ _5064_/A vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6545_ _6545_/A _3268_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3688_ _3688_/A _3688_/B vssd1 vssd1 vccd1 vccd1 _3688_/X sky130_fd_sc_hd__or2_1
X_5427_ _5427_/A _5427_/B vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__xor2_2
XANTENNA__4098__B _4138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5358_ _5358_/A _5358_/B vssd1 vssd1 vccd1 vccd1 _5359_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4309_ _4309_/A _4309_/B vssd1 vssd1 vccd1 vccd1 _4320_/A sky130_fd_sc_hd__xnor2_1
X_5289_ _5289_/A _5289_/B vssd1 vssd1 vccd1 vccd1 _5290_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6505__24 vssd1 vssd1 vccd1 vccd1 _6505__24/HI _6505_/A sky130_fd_sc_hd__conb_1
XFILLER_99_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3905__B _4063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__A _3195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4660_ _4689_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__and2b_1
X_6590__106 vssd1 vssd1 vccd1 vccd1 _6590__106/HI _6590_/A sky130_fd_sc_hd__conb_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ _3611_/A vssd1 vssd1 vccd1 vccd1 _3632_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4591_ _4603_/B _4591_/B vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__xor2_1
X_6330_ _6345_/CLK _6330_/D vssd1 vssd1 vccd1 vccd1 _6330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3542_ _3536_/X _3535_/Y _3534_/Y _3525_/Y vssd1 vssd1 vccd1 vccd1 _3543_/C sky130_fd_sc_hd__o211ai_1
X_3473_ _3473_/A _3473_/B vssd1 vssd1 vccd1 vccd1 _3474_/B sky130_fd_sc_hd__nor2_1
X_6261_ _6267_/A _6261_/B vssd1 vssd1 vccd1 vccd1 _6261_/Y sky130_fd_sc_hd__nor2_1
X_5212_ _5212_/A _5212_/B vssd1 vssd1 vccd1 vccd1 _5242_/B sky130_fd_sc_hd__nor2_1
X_6192_ _6192_/A vssd1 vssd1 vccd1 vccd1 _6353_/D sky130_fd_sc_hd__clkbuf_1
X_5143_ _5136_/A _5142_/Y _4062_/A _5183_/B vssd1 vssd1 vccd1 vccd1 _5151_/A sky130_fd_sc_hd__o211ai_2
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4927__A _5134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5074_ _5074_/A _5074_/B vssd1 vssd1 vccd1 vccd1 _5075_/C sky130_fd_sc_hd__xor2_1
XFILLER_57_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4025_ _5243_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4365__C _4365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5976_ _5974_/X _5976_/B vssd1 vssd1 vccd1 vccd1 _5977_/A sky130_fd_sc_hd__and2b_1
X_4927_ _5134_/B vssd1 vssd1 vccd1 vccd1 _5278_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3278__A _3282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4858_ _4855_/A _4855_/B _4855_/C vssd1 vssd1 vccd1 vccd1 _4858_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3809_ _3810_/A _3810_/B _3810_/C vssd1 vssd1 vccd1 vccd1 _3811_/A sky130_fd_sc_hd__a21oi_1
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4789_ _4815_/A _4787_/X _4788_/X vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__a21boi_1
X_6528_ _6528_/A _3237_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4572__A _5634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_366 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3188__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6577__93 vssd1 vssd1 vccd1 vccd1 _6577__93/HI _6577_/A sky130_fd_sc_hd__conb_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _5813_/X _5747_/X _5749_/Y _5814_/X vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_388 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5761_ _5901_/A _5700_/X _5760_/X _5706_/X vssd1 vssd1 vccd1 vccd1 _5761_/X sky130_fd_sc_hd__o2bb2a_1
X_4712_ _4712_/A _4712_/B vssd1 vssd1 vccd1 vccd1 _4719_/C sky130_fd_sc_hd__nor2_1
X_5692_ _5819_/A vssd1 vssd1 vccd1 vccd1 _5777_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4643_ _4785_/D vssd1 vssd1 vccd1 vccd1 _4692_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4574_ _4574_/A _4574_/B vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__and2_1
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6313_ _6359_/CLK _6313_/D vssd1 vssd1 vccd1 vccd1 _6313_/Q sky130_fd_sc_hd__dfxtp_1
X_3525_ _3527_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _3525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6244_/A vssd1 vssd1 vccd1 vccd1 _6267_/A sky130_fd_sc_hd__clkbuf_2
X_6496__15 vssd1 vssd1 vccd1 vccd1 _6496__15/HI _6496_/A sky130_fd_sc_hd__conb_1
X_3456_ _3386_/A _3391_/A _6299_/Q vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6175_ _6175_/A vssd1 vssd1 vccd1 vccd1 _6347_/D sky130_fd_sc_hd__clkbuf_1
X_3387_ _3387_/A vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5126_ _5125_/A _5125_/B _5125_/C vssd1 vssd1 vccd1 vccd1 _5270_/A sky130_fd_sc_hd__a21o_1
XFILLER_69_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5057_ _5554_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _5082_/A sky130_fd_sc_hd__nand2_1
X_4008_ _4009_/A _4008_/B _4008_/C vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__nand3_1
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5959_ _5959_/A _5959_/B _5959_/C vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__and3_1
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5756__A1 _5710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3310_ _3312_/A vssd1 vssd1 vccd1 vccd1 _3310_/Y sky130_fd_sc_hd__inv_2
X_4290_ _4292_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__and2b_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3245_/A vssd1 vssd1 vccd1 vccd1 _3241_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6596__112 vssd1 vssd1 vccd1 vccd1 _6596__112/HI _6596_/A sky130_fd_sc_hd__conb_1
XFILLER_34_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5813_ _5770_/A _5813_/B _6060_/A vssd1 vssd1 vccd1 vccd1 _5813_/X sky130_fd_sc_hd__and3b_1
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5744_ _6363_/Q _5838_/B _5744_/C vssd1 vssd1 vccd1 vccd1 _5744_/X sky130_fd_sc_hd__or3_1
X_5675_ _5675_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__nor2_1
X_4626_ _4626_/A _5710_/A _5710_/B vssd1 vssd1 vccd1 vccd1 _5757_/A sky130_fd_sc_hd__or3_1
X_4557_ _4978_/A vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__buf_2
XFILLER_104_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4488_ _4488_/A _4488_/B vssd1 vssd1 vccd1 vccd1 _4489_/B sky130_fd_sc_hd__xnor2_2
X_3508_ _3508_/A _3508_/B _3507_/X vssd1 vssd1 vccd1 vccd1 _3508_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3291__A _3294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6227_ _6366_/Q _6365_/Q _6227_/C vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__and3_1
X_3439_ _3549_/C vssd1 vssd1 vccd1 vccd1 _3652_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6334_/Q _6333_/Q _6336_/Q _6335_/Q vssd1 vssd1 vccd1 vccd1 _6158_/X sky130_fd_sc_hd__and4_1
XFILLER_111_190 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5109_ _5109_/A _5109_/B _5109_/C vssd1 vssd1 vccd1 vccd1 _5118_/A sky130_fd_sc_hd__and3_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6089_ _6314_/Q _6189_/B vssd1 vssd1 vccd1 vccd1 _6090_/A sky130_fd_sc_hd__and2_1
XFILLER_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5011__A _5011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3461__A2 _4814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4850__A _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6547__63 vssd1 vssd1 vccd1 vccd1 _6547__63/HI _6547_/A sky130_fd_sc_hd__conb_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5681__A _5737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3790_ _5011_/A _4235_/B _3947_/B _5007_/A vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__a22o_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5294__C _5505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5460_ _5462_/A _5462_/B _5459_/X vssd1 vssd1 vccd1 vccd1 _5533_/B sky130_fd_sc_hd__a21boi_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4411_ _4411_/A _4435_/A vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__xor2_1
X_5391_ _5394_/A _5440_/B vssd1 vssd1 vccd1 vccd1 _5393_/A sky130_fd_sc_hd__nand2_1
X_4342_ _4409_/B vssd1 vssd1 vccd1 vccd1 _4580_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4273_ _4273_/A _4273_/B vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__xor2_2
XFILLER_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3224_ _3226_/A vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6012_ _6057_/A _6012_/B vssd1 vssd1 vccd1 vccd1 _6012_/Y sky130_fd_sc_hd__nand2_1
.ends

